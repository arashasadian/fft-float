library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


package fftpackage is
    constant PI : integer := 180;
    constant TwoPI : integer := 360;
    constant ROWS, COLS : integer := 512;
    constant STEP : integer := 9;
    -- constant THRESHOLD : float32 := to_float(100);
    constant bitWidth : integer := 26;
    --type array_of_float32 is array(natural range <>) of float32;
    type array_of_slv is array (natural range <>) of std_logic_vector(bitWidth-1 downto 0);
    type array_2d_slv is array (natural range <>) of array_of_slv;
    type array_of_integer is array(natural range <>) of integer;
    -- type array_2d_float is array(natural range <>) of array_of_float32;
    type fft_state is (RESET_STATE, IDLE, INIT, INIT2, BUSY1, BUSY2);
    type fft2d_state is (IDLE, TRANSPOSE ,FFT1_RESET, FAKE1, FFT1, FFT1_P, TRANSPOSE1, FFT2_RESET,FAKE, FFT2, FFT2_P);
    
    component transpose_matrix is
      generic ( ROWS : integer ; COLS : integer );
    port (
      enable : in std_logic;
      buffer_real_in  : in array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
      buffer_imag_in  : in array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
      buffer_real_out : out array_2d_slv(COLS-1 downto 0)(ROWS-1 downto 0);
      buffer_imag_out : out array_2d_slv(COLS-1 downto 0)(ROWS-1 downto 0)
    ) ;
    end component transpose_matrix;

    -- component filter is
    --   generic ( ROWS : integer ; COLS : integer );
    --   port (
    --     enable : in std_logic;
    --     buffer_real_in  : in array_2d_float(ROWS-1 downto 0)(COLS-1 downto 0);
    --     buffer_imag_in  : in array_2d_float(ROWS-1 downto 0)(COLS-1 downto 0);
    --     buffer_real_out : out array_2d_float(COLS-1 downto 0)(ROWS-1 downto 0);
    --     buffer_imag_out : out array_2d_float(COLS-1 downto 0)(ROWS-1 downto 0)
    --   ) ;
    -- end component filter;

    component butterfly is
      generic(bitWidth : integer := 32);
      port (
        clk : in std_logic;
        input1_real : in std_logic_vector(bitWidth-1 downto 0);
        input1_imag : in std_logic_vector(bitWidth-1 downto 0);
        input2_real : in std_logic_vector(bitWidth-1 downto 0);
        input2_imag : in std_logic_vector(bitWidth-1 downto 0);
        coefficient_real : in std_logic_vector(bitWidth-1 downto 0);
        coefficient_imag : in std_logic_vector(bitWidth-1 downto 0);
        output1_real : out std_logic_vector(bitWidth-1 downto 0);
        output1_imag : out std_logic_vector(bitWidth-1 downto 0);
        output2_real : out std_logic_vector(bitWidth-1 downto 0);
        output2_imag : out std_logic_vector(bitWidth-1 downto 0)
      ) ;
    end component butterfly;

      component fft is
        generic ( N : integer := 8; step : integer := 3);
        port (
          clk : in std_logic;
          reset : in std_logic;
          input_array_real : in array_of_slv(N - 1 downto 0);
          input_array_imag : in array_of_slv(N - 1 downto 0);
          output_array_real : out array_of_slv(N - 1 downto 0);
          output_array_imag : out array_of_slv(N - 1 downto 0);
          done : out std_logic
        ) ;
      end component fft;

      component fft_top is
      generic ( ROWS : integer; COLS : integer);
      port (
        clk : in std_logic;
        reset : in std_logic;
        enable : in std_logic;
        buffer_real_in  : in array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
        buffer_imag_in  : in array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
        buffer_real_out : out array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
        buffer_imag_out : out array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
        done : out std_logic
      );
    end component fft_top;

  component ifft2d is
    generic ( ROWS : integer ; COLS : integer );
    port (
      clk : in std_logic;
      reset : in std_logic;
      enable : in std_logic;
      input_array_real : in array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
      input_array_imag : in array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
      output_array_real : out array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
      output_array_imag : out array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
      done : out std_logic
    ) ;
  end component ifft2d;


    component ifft is
      generic ( N : integer := 8; step : integer := 3);
      port (
        clk : in std_logic;
        reset : in std_logic;
        input_array_real : in array_of_slv(N - 1 downto 0);
        input_array_imag : in array_of_slv(N - 1 downto 0);
        output_array_real : out array_of_slv(N - 1 downto 0);
        output_array_imag : out array_of_slv(N - 1 downto 0);
        done : out std_logic
      ) ;
    end component ifft;

    component ifft_top is
      generic ( ROWS : integer; COLS : integer);
      port (
        clk : in std_logic;
        reset : in std_logic;
        enable : in std_logic;
        buffer_real_in  : in array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
        buffer_imag_in  : in array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
        buffer_real_out : out array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
        buffer_imag_out : out array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
        done : out std_logic
      ) ;
      end component ifft_top;

    component fft2d is
      generic ( ROWS : integer ; COLS : integer );
      port (
      clk : in std_logic;
      reset : in std_logic;
      enable : in std_logic;
      input_array_real : in array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
      input_array_imag : in array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
      output_array_real : out array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
      output_array_imag : out array_2d_slv(ROWS-1 downto 0)(COLS-1 downto 0);
      done : out std_logic
    ) ;
    end component fft2d;
    -- signal middle_index_rom : array_of_integer(7 downto 0);
    -- signal output_index_rom : array_of_integer(7 downto 0);
    -- signal input_index_rom : array_of_integer(7 downto 0);
    signal sin_rom, cos_rom : array_of_slv(360 downto 0);
    -- signal buffer_2d_real, buffer_2d_imag : array_2d_float(ROWS-1 downto 0)(COLS-1 downto 0);
    procedure trigonometrics_rom_generator (
      signal enable : in std_logic ;
      signal s_rom, c_rom : inout array_of_slv(360 downto 0));   
      -- procedure buffer_init(reset : in std_logic; signal re, im : inout array_2d_float(ROWS-1 downto 0)(COLS-1 downto 0));

end package fftpackage;

package body fftpackage is 
  
  -- procedure buffer_init(reset : in std_logic; signal re, im : inout array_2d_float(ROWS-1 downto 0)(COLS-1 downto 0))
  --     is begin
  --       for i in 0 to ROWS-1 loop
  --         for j in 0 to COLS -1 loop
  --             re(i)(j) <= to_float(i * j);
  --             im(i)(j) <= to_float(i - j);
  --             report "i = " & integer'image(i);
  --             report "j = " & integer'image(j);
  --         end loop;
  --     end loop;
  -- end procedure;


  procedure trigonometrics_rom_generator (
      signal enable : in std_logic ;
      signal s_rom, c_rom : inout array_of_slv(360 downto 0)
      )is
    begin
      if rising_edge(enable) then 
      s_rom(0) <= std_logic_vector(to_signed(0,bitWidth));
      s_rom(1) <= std_logic_vector(to_signed(4,bitWidth));
      s_rom(2) <= std_logic_vector(to_signed(8,bitWidth));
      s_rom(3) <= std_logic_vector(to_signed(13,bitWidth));
      s_rom(4) <= std_logic_vector(to_signed(17,bitWidth));
      s_rom(5) <= std_logic_vector(to_signed(22,bitWidth));
      s_rom(6) <= std_logic_vector(to_signed(26,bitWidth));
      s_rom(7) <= std_logic_vector(to_signed(31,bitWidth));
      s_rom(8) <= std_logic_vector(to_signed(35,bitWidth));
      s_rom(9) <= std_logic_vector(to_signed(39,bitWidth));
      s_rom(10) <= std_logic_vector(to_signed(44,bitWidth));
      s_rom(11) <= std_logic_vector(to_signed(48,bitWidth));
      s_rom(12) <= std_logic_vector(to_signed(53,bitWidth));
      s_rom(13) <= std_logic_vector(to_signed(57,bitWidth));
      s_rom(14) <= std_logic_vector(to_signed(61,bitWidth));
      s_rom(15) <= std_logic_vector(to_signed(65,bitWidth));
      s_rom(16) <= std_logic_vector(to_signed(70,bitWidth));
      s_rom(17) <= std_logic_vector(to_signed(74,bitWidth));
      s_rom(18) <= std_logic_vector(to_signed(78,bitWidth));
      s_rom(19) <= std_logic_vector(to_signed(83,bitWidth));
      s_rom(20) <= std_logic_vector(to_signed(87,bitWidth));
      s_rom(21) <= std_logic_vector(to_signed(91,bitWidth));
      s_rom(22) <= std_logic_vector(to_signed(95,bitWidth));
      s_rom(23) <= std_logic_vector(to_signed(99,bitWidth));
      s_rom(24) <= std_logic_vector(to_signed(103,bitWidth));
      s_rom(25) <= std_logic_vector(to_signed(107,bitWidth));
      s_rom(26) <= std_logic_vector(to_signed(111,bitWidth));
      s_rom(27) <= std_logic_vector(to_signed(115,bitWidth));
      s_rom(28) <= std_logic_vector(to_signed(119,bitWidth));
      s_rom(29) <= std_logic_vector(to_signed(123,bitWidth));
      s_rom(30) <= std_logic_vector(to_signed(127,bitWidth));
      s_rom(31) <= std_logic_vector(to_signed(131,bitWidth));
      s_rom(32) <= std_logic_vector(to_signed(135,bitWidth));
      s_rom(33) <= std_logic_vector(to_signed(138,bitWidth));
      s_rom(34) <= std_logic_vector(to_signed(142,bitWidth));
      s_rom(35) <= std_logic_vector(to_signed(146,bitWidth));
      s_rom(36) <= std_logic_vector(to_signed(149,bitWidth));
      s_rom(37) <= std_logic_vector(to_signed(153,bitWidth));
      s_rom(38) <= std_logic_vector(to_signed(156,bitWidth));
      s_rom(39) <= std_logic_vector(to_signed(160,bitWidth));
      s_rom(40) <= std_logic_vector(to_signed(163,bitWidth));
      s_rom(41) <= std_logic_vector(to_signed(167,bitWidth));
      s_rom(42) <= std_logic_vector(to_signed(170,bitWidth));
      s_rom(43) <= std_logic_vector(to_signed(173,bitWidth));
      s_rom(44) <= std_logic_vector(to_signed(177,bitWidth));
      s_rom(45) <= std_logic_vector(to_signed(180,bitWidth));
      s_rom(46) <= std_logic_vector(to_signed(183,bitWidth));
      s_rom(47) <= std_logic_vector(to_signed(186,bitWidth));
      s_rom(48) <= std_logic_vector(to_signed(189,bitWidth));
      s_rom(49) <= std_logic_vector(to_signed(192,bitWidth));
      s_rom(50) <= std_logic_vector(to_signed(195,bitWidth));
      s_rom(51) <= std_logic_vector(to_signed(198,bitWidth));
      s_rom(52) <= std_logic_vector(to_signed(200,bitWidth));
      s_rom(53) <= std_logic_vector(to_signed(203,bitWidth));
      s_rom(54) <= std_logic_vector(to_signed(206,bitWidth));
      s_rom(55) <= std_logic_vector(to_signed(208,bitWidth));
      s_rom(56) <= std_logic_vector(to_signed(211,bitWidth));
      s_rom(57) <= std_logic_vector(to_signed(213,bitWidth));
      s_rom(58) <= std_logic_vector(to_signed(216,bitWidth));
      s_rom(59) <= std_logic_vector(to_signed(218,bitWidth));
      s_rom(60) <= std_logic_vector(to_signed(220,bitWidth));
      s_rom(61) <= std_logic_vector(to_signed(223,bitWidth));
      s_rom(62) <= std_logic_vector(to_signed(225,bitWidth));
      s_rom(63) <= std_logic_vector(to_signed(227,bitWidth));
      s_rom(64) <= std_logic_vector(to_signed(229,bitWidth));
      s_rom(65) <= std_logic_vector(to_signed(231,bitWidth));
      s_rom(66) <= std_logic_vector(to_signed(232,bitWidth));
      s_rom(67) <= std_logic_vector(to_signed(234,bitWidth));
      s_rom(68) <= std_logic_vector(to_signed(236,bitWidth));
      s_rom(69) <= std_logic_vector(to_signed(238,bitWidth));
      s_rom(70) <= std_logic_vector(to_signed(239,bitWidth));
      s_rom(71) <= std_logic_vector(to_signed(241,bitWidth));
      s_rom(72) <= std_logic_vector(to_signed(242,bitWidth));
      s_rom(73) <= std_logic_vector(to_signed(243,bitWidth));
      s_rom(74) <= std_logic_vector(to_signed(245,bitWidth));
      s_rom(75) <= std_logic_vector(to_signed(246,bitWidth));
      s_rom(76) <= std_logic_vector(to_signed(247,bitWidth));
      s_rom(77) <= std_logic_vector(to_signed(248,bitWidth));
      s_rom(78) <= std_logic_vector(to_signed(249,bitWidth));
      s_rom(79) <= std_logic_vector(to_signed(250,bitWidth));
      s_rom(80) <= std_logic_vector(to_signed(251,bitWidth));
      s_rom(81) <= std_logic_vector(to_signed(251,bitWidth));
      s_rom(82) <= std_logic_vector(to_signed(252,bitWidth));
      s_rom(83) <= std_logic_vector(to_signed(253,bitWidth));
      s_rom(84) <= std_logic_vector(to_signed(253,bitWidth));
      s_rom(85) <= std_logic_vector(to_signed(254,bitWidth));
      s_rom(86) <= std_logic_vector(to_signed(254,bitWidth));
      s_rom(87) <= std_logic_vector(to_signed(254,bitWidth));
      s_rom(88) <= std_logic_vector(to_signed(254,bitWidth));
      s_rom(89) <= std_logic_vector(to_signed(254,bitWidth));
      s_rom(90) <= std_logic_vector(to_signed(255,bitWidth));
      s_rom(91) <= std_logic_vector(to_signed(254,bitWidth));
      s_rom(92) <= std_logic_vector(to_signed(254,bitWidth));
      s_rom(93) <= std_logic_vector(to_signed(254,bitWidth));
      s_rom(94) <= std_logic_vector(to_signed(254,bitWidth));
      s_rom(95) <= std_logic_vector(to_signed(254,bitWidth));
      s_rom(96) <= std_logic_vector(to_signed(253,bitWidth));
      s_rom(97) <= std_logic_vector(to_signed(253,bitWidth));
      s_rom(98) <= std_logic_vector(to_signed(252,bitWidth));
      s_rom(99) <= std_logic_vector(to_signed(251,bitWidth));
      s_rom(100) <= std_logic_vector(to_signed(251,bitWidth));
      s_rom(101) <= std_logic_vector(to_signed(250,bitWidth));
      s_rom(102) <= std_logic_vector(to_signed(249,bitWidth));
      s_rom(103) <= std_logic_vector(to_signed(248,bitWidth));
      s_rom(104) <= std_logic_vector(to_signed(247,bitWidth));
      s_rom(105) <= std_logic_vector(to_signed(246,bitWidth));
      s_rom(106) <= std_logic_vector(to_signed(245,bitWidth));
      s_rom(107) <= std_logic_vector(to_signed(243,bitWidth));
      s_rom(108) <= std_logic_vector(to_signed(242,bitWidth));
      s_rom(109) <= std_logic_vector(to_signed(241,bitWidth));
      s_rom(110) <= std_logic_vector(to_signed(239,bitWidth));
      s_rom(111) <= std_logic_vector(to_signed(238,bitWidth));
      s_rom(112) <= std_logic_vector(to_signed(236,bitWidth));
      s_rom(113) <= std_logic_vector(to_signed(234,bitWidth));
      s_rom(114) <= std_logic_vector(to_signed(232,bitWidth));
      s_rom(115) <= std_logic_vector(to_signed(231,bitWidth));
      s_rom(116) <= std_logic_vector(to_signed(229,bitWidth));
      s_rom(117) <= std_logic_vector(to_signed(227,bitWidth));
      s_rom(118) <= std_logic_vector(to_signed(225,bitWidth));
      s_rom(119) <= std_logic_vector(to_signed(223,bitWidth));
      s_rom(120) <= std_logic_vector(to_signed(220,bitWidth));
      s_rom(121) <= std_logic_vector(to_signed(218,bitWidth));
      s_rom(122) <= std_logic_vector(to_signed(216,bitWidth));
      s_rom(123) <= std_logic_vector(to_signed(213,bitWidth));
      s_rom(124) <= std_logic_vector(to_signed(211,bitWidth));
      s_rom(125) <= std_logic_vector(to_signed(208,bitWidth));
      s_rom(126) <= std_logic_vector(to_signed(206,bitWidth));
      s_rom(127) <= std_logic_vector(to_signed(203,bitWidth));
      s_rom(128) <= std_logic_vector(to_signed(200,bitWidth));
      s_rom(129) <= std_logic_vector(to_signed(198,bitWidth));
      s_rom(130) <= std_logic_vector(to_signed(195,bitWidth));
      s_rom(131) <= std_logic_vector(to_signed(192,bitWidth));
      s_rom(132) <= std_logic_vector(to_signed(189,bitWidth));
      s_rom(133) <= std_logic_vector(to_signed(186,bitWidth));
      s_rom(134) <= std_logic_vector(to_signed(183,bitWidth));
      s_rom(135) <= std_logic_vector(to_signed(180,bitWidth));
      s_rom(136) <= std_logic_vector(to_signed(177,bitWidth));
      s_rom(137) <= std_logic_vector(to_signed(173,bitWidth));
      s_rom(138) <= std_logic_vector(to_signed(170,bitWidth));
      s_rom(139) <= std_logic_vector(to_signed(167,bitWidth));
      s_rom(140) <= std_logic_vector(to_signed(163,bitWidth));
      s_rom(141) <= std_logic_vector(to_signed(160,bitWidth));
      s_rom(142) <= std_logic_vector(to_signed(156,bitWidth));
      s_rom(143) <= std_logic_vector(to_signed(153,bitWidth));
      s_rom(144) <= std_logic_vector(to_signed(149,bitWidth));
      s_rom(145) <= std_logic_vector(to_signed(146,bitWidth));
      s_rom(146) <= std_logic_vector(to_signed(142,bitWidth));
      s_rom(147) <= std_logic_vector(to_signed(138,bitWidth));
      s_rom(148) <= std_logic_vector(to_signed(135,bitWidth));
      s_rom(149) <= std_logic_vector(to_signed(131,bitWidth));
      s_rom(150) <= std_logic_vector(to_signed(127,bitWidth));
      s_rom(151) <= std_logic_vector(to_signed(123,bitWidth));
      s_rom(152) <= std_logic_vector(to_signed(119,bitWidth));
      s_rom(153) <= std_logic_vector(to_signed(115,bitWidth));
      s_rom(154) <= std_logic_vector(to_signed(111,bitWidth));
      s_rom(155) <= std_logic_vector(to_signed(107,bitWidth));
      s_rom(156) <= std_logic_vector(to_signed(103,bitWidth));
      s_rom(157) <= std_logic_vector(to_signed(99,bitWidth));
      s_rom(158) <= std_logic_vector(to_signed(95,bitWidth));
      s_rom(159) <= std_logic_vector(to_signed(91,bitWidth));
      s_rom(160) <= std_logic_vector(to_signed(87,bitWidth));
      s_rom(161) <= std_logic_vector(to_signed(83,bitWidth));
      s_rom(162) <= std_logic_vector(to_signed(78,bitWidth));
      s_rom(163) <= std_logic_vector(to_signed(74,bitWidth));
      s_rom(164) <= std_logic_vector(to_signed(70,bitWidth));
      s_rom(165) <= std_logic_vector(to_signed(65,bitWidth));
      s_rom(166) <= std_logic_vector(to_signed(61,bitWidth));
      s_rom(167) <= std_logic_vector(to_signed(57,bitWidth));
      s_rom(168) <= std_logic_vector(to_signed(53,bitWidth));
      s_rom(169) <= std_logic_vector(to_signed(48,bitWidth));
      s_rom(170) <= std_logic_vector(to_signed(44,bitWidth));
      s_rom(171) <= std_logic_vector(to_signed(39,bitWidth));
      s_rom(172) <= std_logic_vector(to_signed(35,bitWidth));
      s_rom(173) <= std_logic_vector(to_signed(31,bitWidth));
      s_rom(174) <= std_logic_vector(to_signed(26,bitWidth));
      s_rom(175) <= std_logic_vector(to_signed(22,bitWidth));
      s_rom(176) <= std_logic_vector(to_signed(17,bitWidth));
      s_rom(177) <= std_logic_vector(to_signed(13,bitWidth));
      s_rom(178) <= std_logic_vector(to_signed(8,bitWidth));
      s_rom(179) <= std_logic_vector(to_signed(4,bitWidth));
      s_rom(180) <= std_logic_vector(to_signed(0,bitWidth));
      s_rom(181) <= std_logic_vector(to_signed(-4,bitWidth));
      s_rom(182) <= std_logic_vector(to_signed(-8,bitWidth));
      s_rom(183) <= std_logic_vector(to_signed(-13,bitWidth));
      s_rom(184) <= std_logic_vector(to_signed(-17,bitWidth));
      s_rom(185) <= std_logic_vector(to_signed(-22,bitWidth));
      s_rom(186) <= std_logic_vector(to_signed(-26,bitWidth));
      s_rom(187) <= std_logic_vector(to_signed(-31,bitWidth));
      s_rom(188) <= std_logic_vector(to_signed(-35,bitWidth));
      s_rom(189) <= std_logic_vector(to_signed(-39,bitWidth));
      s_rom(190) <= std_logic_vector(to_signed(-44,bitWidth));
      s_rom(191) <= std_logic_vector(to_signed(-48,bitWidth));
      s_rom(192) <= std_logic_vector(to_signed(-53,bitWidth));
      s_rom(193) <= std_logic_vector(to_signed(-57,bitWidth));
      s_rom(194) <= std_logic_vector(to_signed(-61,bitWidth));
      s_rom(195) <= std_logic_vector(to_signed(-65,bitWidth));
      s_rom(196) <= std_logic_vector(to_signed(-70,bitWidth));
      s_rom(197) <= std_logic_vector(to_signed(-74,bitWidth));
      s_rom(198) <= std_logic_vector(to_signed(-78,bitWidth));
      s_rom(199) <= std_logic_vector(to_signed(-83,bitWidth));
      s_rom(200) <= std_logic_vector(to_signed(-87,bitWidth));
      s_rom(201) <= std_logic_vector(to_signed(-91,bitWidth));
      s_rom(202) <= std_logic_vector(to_signed(-95,bitWidth));
      s_rom(203) <= std_logic_vector(to_signed(-99,bitWidth));
      s_rom(204) <= std_logic_vector(to_signed(-103,bitWidth));
      s_rom(205) <= std_logic_vector(to_signed(-107,bitWidth));
      s_rom(206) <= std_logic_vector(to_signed(-111,bitWidth));
      s_rom(207) <= std_logic_vector(to_signed(-115,bitWidth));
      s_rom(208) <= std_logic_vector(to_signed(-119,bitWidth));
      s_rom(209) <= std_logic_vector(to_signed(-123,bitWidth));
      s_rom(210) <= std_logic_vector(to_signed(-127,bitWidth));
      s_rom(211) <= std_logic_vector(to_signed(-131,bitWidth));
      s_rom(212) <= std_logic_vector(to_signed(-135,bitWidth));
      s_rom(213) <= std_logic_vector(to_signed(-138,bitWidth));
      s_rom(214) <= std_logic_vector(to_signed(-142,bitWidth));
      s_rom(215) <= std_logic_vector(to_signed(-146,bitWidth));
      s_rom(216) <= std_logic_vector(to_signed(-149,bitWidth));
      s_rom(217) <= std_logic_vector(to_signed(-153,bitWidth));
      s_rom(218) <= std_logic_vector(to_signed(-156,bitWidth));
      s_rom(219) <= std_logic_vector(to_signed(-160,bitWidth));
      s_rom(220) <= std_logic_vector(to_signed(-163,bitWidth));
      s_rom(221) <= std_logic_vector(to_signed(-167,bitWidth));
      s_rom(222) <= std_logic_vector(to_signed(-170,bitWidth));
      s_rom(223) <= std_logic_vector(to_signed(-173,bitWidth));
      s_rom(224) <= std_logic_vector(to_signed(-177,bitWidth));
      s_rom(225) <= std_logic_vector(to_signed(-180,bitWidth));
      s_rom(226) <= std_logic_vector(to_signed(-183,bitWidth));
      s_rom(227) <= std_logic_vector(to_signed(-186,bitWidth));
      s_rom(228) <= std_logic_vector(to_signed(-189,bitWidth));
      s_rom(229) <= std_logic_vector(to_signed(-192,bitWidth));
      s_rom(230) <= std_logic_vector(to_signed(-195,bitWidth));
      s_rom(231) <= std_logic_vector(to_signed(-198,bitWidth));
      s_rom(232) <= std_logic_vector(to_signed(-200,bitWidth));
      s_rom(233) <= std_logic_vector(to_signed(-203,bitWidth));
      s_rom(234) <= std_logic_vector(to_signed(-206,bitWidth));
      s_rom(235) <= std_logic_vector(to_signed(-208,bitWidth));
      s_rom(236) <= std_logic_vector(to_signed(-211,bitWidth));
      s_rom(237) <= std_logic_vector(to_signed(-213,bitWidth));
      s_rom(238) <= std_logic_vector(to_signed(-216,bitWidth));
      s_rom(239) <= std_logic_vector(to_signed(-218,bitWidth));
      s_rom(240) <= std_logic_vector(to_signed(-220,bitWidth));
      s_rom(241) <= std_logic_vector(to_signed(-223,bitWidth));
      s_rom(242) <= std_logic_vector(to_signed(-225,bitWidth));
      s_rom(243) <= std_logic_vector(to_signed(-227,bitWidth));
      s_rom(244) <= std_logic_vector(to_signed(-229,bitWidth));
      s_rom(245) <= std_logic_vector(to_signed(-231,bitWidth));
      s_rom(246) <= std_logic_vector(to_signed(-232,bitWidth));
      s_rom(247) <= std_logic_vector(to_signed(-234,bitWidth));
      s_rom(248) <= std_logic_vector(to_signed(-236,bitWidth));
      s_rom(249) <= std_logic_vector(to_signed(-238,bitWidth));
      s_rom(250) <= std_logic_vector(to_signed(-239,bitWidth));
      s_rom(251) <= std_logic_vector(to_signed(-241,bitWidth));
      s_rom(252) <= std_logic_vector(to_signed(-242,bitWidth));
      s_rom(253) <= std_logic_vector(to_signed(-243,bitWidth));
      s_rom(254) <= std_logic_vector(to_signed(-245,bitWidth));
      s_rom(255) <= std_logic_vector(to_signed(-246,bitWidth));
      s_rom(256) <= std_logic_vector(to_signed(-247,bitWidth));
      s_rom(257) <= std_logic_vector(to_signed(-248,bitWidth));
      s_rom(258) <= std_logic_vector(to_signed(-249,bitWidth));
      s_rom(259) <= std_logic_vector(to_signed(-250,bitWidth));
      s_rom(260) <= std_logic_vector(to_signed(-251,bitWidth));
      s_rom(261) <= std_logic_vector(to_signed(-251,bitWidth));
      s_rom(262) <= std_logic_vector(to_signed(-252,bitWidth));
      s_rom(263) <= std_logic_vector(to_signed(-253,bitWidth));
      s_rom(264) <= std_logic_vector(to_signed(-253,bitWidth));
      s_rom(265) <= std_logic_vector(to_signed(-254,bitWidth));
      s_rom(266) <= std_logic_vector(to_signed(-254,bitWidth));
      s_rom(267) <= std_logic_vector(to_signed(-254,bitWidth));
      s_rom(268) <= std_logic_vector(to_signed(-254,bitWidth));
      s_rom(269) <= std_logic_vector(to_signed(-254,bitWidth));
      s_rom(270) <= std_logic_vector(to_signed(-255,bitWidth));
      s_rom(271) <= std_logic_vector(to_signed(-254,bitWidth));
      s_rom(272) <= std_logic_vector(to_signed(-254,bitWidth));
      s_rom(273) <= std_logic_vector(to_signed(-254,bitWidth));
      s_rom(274) <= std_logic_vector(to_signed(-254,bitWidth));
      s_rom(275) <= std_logic_vector(to_signed(-254,bitWidth));
      s_rom(276) <= std_logic_vector(to_signed(-253,bitWidth));
      s_rom(277) <= std_logic_vector(to_signed(-253,bitWidth));
      s_rom(278) <= std_logic_vector(to_signed(-252,bitWidth));
      s_rom(279) <= std_logic_vector(to_signed(-251,bitWidth));
      s_rom(280) <= std_logic_vector(to_signed(-251,bitWidth));
      s_rom(281) <= std_logic_vector(to_signed(-250,bitWidth));
      s_rom(282) <= std_logic_vector(to_signed(-249,bitWidth));
      s_rom(283) <= std_logic_vector(to_signed(-248,bitWidth));
      s_rom(284) <= std_logic_vector(to_signed(-247,bitWidth));
      s_rom(285) <= std_logic_vector(to_signed(-246,bitWidth));
      s_rom(286) <= std_logic_vector(to_signed(-245,bitWidth));
      s_rom(287) <= std_logic_vector(to_signed(-243,bitWidth));
      s_rom(288) <= std_logic_vector(to_signed(-242,bitWidth));
      s_rom(289) <= std_logic_vector(to_signed(-241,bitWidth));
      s_rom(290) <= std_logic_vector(to_signed(-239,bitWidth));
      s_rom(291) <= std_logic_vector(to_signed(-238,bitWidth));
      s_rom(292) <= std_logic_vector(to_signed(-236,bitWidth));
      s_rom(293) <= std_logic_vector(to_signed(-234,bitWidth));
      s_rom(294) <= std_logic_vector(to_signed(-232,bitWidth));
      s_rom(295) <= std_logic_vector(to_signed(-231,bitWidth));
      s_rom(296) <= std_logic_vector(to_signed(-229,bitWidth));
      s_rom(297) <= std_logic_vector(to_signed(-227,bitWidth));
      s_rom(298) <= std_logic_vector(to_signed(-225,bitWidth));
      s_rom(299) <= std_logic_vector(to_signed(-223,bitWidth));
      s_rom(300) <= std_logic_vector(to_signed(-220,bitWidth));
      s_rom(301) <= std_logic_vector(to_signed(-218,bitWidth));
      s_rom(302) <= std_logic_vector(to_signed(-216,bitWidth));
      s_rom(303) <= std_logic_vector(to_signed(-213,bitWidth));
      s_rom(304) <= std_logic_vector(to_signed(-211,bitWidth));
      s_rom(305) <= std_logic_vector(to_signed(-208,bitWidth));
      s_rom(306) <= std_logic_vector(to_signed(-206,bitWidth));
      s_rom(307) <= std_logic_vector(to_signed(-203,bitWidth));
      s_rom(308) <= std_logic_vector(to_signed(-200,bitWidth));
      s_rom(309) <= std_logic_vector(to_signed(-198,bitWidth));
      s_rom(310) <= std_logic_vector(to_signed(-195,bitWidth));
      s_rom(311) <= std_logic_vector(to_signed(-192,bitWidth));
      s_rom(312) <= std_logic_vector(to_signed(-189,bitWidth));
      s_rom(313) <= std_logic_vector(to_signed(-186,bitWidth));
      s_rom(314) <= std_logic_vector(to_signed(-183,bitWidth));
      s_rom(315) <= std_logic_vector(to_signed(-180,bitWidth));
      s_rom(316) <= std_logic_vector(to_signed(-177,bitWidth));
      s_rom(317) <= std_logic_vector(to_signed(-173,bitWidth));
      s_rom(318) <= std_logic_vector(to_signed(-170,bitWidth));
      s_rom(319) <= std_logic_vector(to_signed(-167,bitWidth));
      s_rom(320) <= std_logic_vector(to_signed(-163,bitWidth));
      s_rom(321) <= std_logic_vector(to_signed(-160,bitWidth));
      s_rom(322) <= std_logic_vector(to_signed(-156,bitWidth));
      s_rom(323) <= std_logic_vector(to_signed(-153,bitWidth));
      s_rom(324) <= std_logic_vector(to_signed(-149,bitWidth));
      s_rom(325) <= std_logic_vector(to_signed(-146,bitWidth));
      s_rom(326) <= std_logic_vector(to_signed(-142,bitWidth));
      s_rom(327) <= std_logic_vector(to_signed(-138,bitWidth));
      s_rom(328) <= std_logic_vector(to_signed(-135,bitWidth));
      s_rom(329) <= std_logic_vector(to_signed(-131,bitWidth));
      s_rom(330) <= std_logic_vector(to_signed(-127,bitWidth));
      s_rom(331) <= std_logic_vector(to_signed(-123,bitWidth));
      s_rom(332) <= std_logic_vector(to_signed(-119,bitWidth));
      s_rom(333) <= std_logic_vector(to_signed(-115,bitWidth));
      s_rom(334) <= std_logic_vector(to_signed(-111,bitWidth));
      s_rom(335) <= std_logic_vector(to_signed(-107,bitWidth));
      s_rom(336) <= std_logic_vector(to_signed(-103,bitWidth));
      s_rom(337) <= std_logic_vector(to_signed(-99,bitWidth));
      s_rom(338) <= std_logic_vector(to_signed(-95,bitWidth));
      s_rom(339) <= std_logic_vector(to_signed(-91,bitWidth));
      s_rom(340) <= std_logic_vector(to_signed(-87,bitWidth));
      s_rom(341) <= std_logic_vector(to_signed(-83,bitWidth));
      s_rom(342) <= std_logic_vector(to_signed(-78,bitWidth));
      s_rom(343) <= std_logic_vector(to_signed(-74,bitWidth));
      s_rom(344) <= std_logic_vector(to_signed(-70,bitWidth));
      s_rom(345) <= std_logic_vector(to_signed(-65,bitWidth));
      s_rom(346) <= std_logic_vector(to_signed(-61,bitWidth));
      s_rom(347) <= std_logic_vector(to_signed(-57,bitWidth));
      s_rom(348) <= std_logic_vector(to_signed(-53,bitWidth));
      s_rom(349) <= std_logic_vector(to_signed(-48,bitWidth));
      s_rom(350) <= std_logic_vector(to_signed(-44,bitWidth));
      s_rom(351) <= std_logic_vector(to_signed(-39,bitWidth));
      s_rom(352) <= std_logic_vector(to_signed(-35,bitWidth));
      s_rom(353) <= std_logic_vector(to_signed(-31,bitWidth));
      s_rom(354) <= std_logic_vector(to_signed(-26,bitWidth));
      s_rom(355) <= std_logic_vector(to_signed(-22,bitWidth));
      s_rom(356) <= std_logic_vector(to_signed(-17,bitWidth));
      s_rom(357) <= std_logic_vector(to_signed(-13,bitWidth));
      s_rom(358) <= std_logic_vector(to_signed(-8,bitWidth));
      s_rom(359) <= std_logic_vector(to_signed(-4,bitWidth));
      s_rom(360) <= std_logic_vector(to_signed(0,bitWidth));

      c_rom(0) <= std_logic_vector(to_signed(255,bitWidth));
      c_rom(1) <= std_logic_vector(to_signed(254,bitWidth));
      c_rom(2) <= std_logic_vector(to_signed(254,bitWidth));
      c_rom(3) <= std_logic_vector(to_signed(254,bitWidth));
      c_rom(4) <= std_logic_vector(to_signed(254,bitWidth));
      c_rom(5) <= std_logic_vector(to_signed(254,bitWidth));
      c_rom(6) <= std_logic_vector(to_signed(253,bitWidth));
      c_rom(7) <= std_logic_vector(to_signed(253,bitWidth));
      c_rom(8) <= std_logic_vector(to_signed(252,bitWidth));
      c_rom(9) <= std_logic_vector(to_signed(251,bitWidth));
      c_rom(10) <= std_logic_vector(to_signed(251,bitWidth));
      c_rom(11) <= std_logic_vector(to_signed(250,bitWidth));
      c_rom(12) <= std_logic_vector(to_signed(249,bitWidth));
      c_rom(13) <= std_logic_vector(to_signed(248,bitWidth));
      c_rom(14) <= std_logic_vector(to_signed(247,bitWidth));
      c_rom(15) <= std_logic_vector(to_signed(246,bitWidth));
      c_rom(16) <= std_logic_vector(to_signed(245,bitWidth));
      c_rom(17) <= std_logic_vector(to_signed(243,bitWidth));
      c_rom(18) <= std_logic_vector(to_signed(242,bitWidth));
      c_rom(19) <= std_logic_vector(to_signed(241,bitWidth));
      c_rom(20) <= std_logic_vector(to_signed(239,bitWidth));
      c_rom(21) <= std_logic_vector(to_signed(238,bitWidth));
      c_rom(22) <= std_logic_vector(to_signed(236,bitWidth));
      c_rom(23) <= std_logic_vector(to_signed(234,bitWidth));
      c_rom(24) <= std_logic_vector(to_signed(232,bitWidth));
      c_rom(25) <= std_logic_vector(to_signed(231,bitWidth));
      c_rom(26) <= std_logic_vector(to_signed(229,bitWidth));
      c_rom(27) <= std_logic_vector(to_signed(227,bitWidth));
      c_rom(28) <= std_logic_vector(to_signed(225,bitWidth));
      c_rom(29) <= std_logic_vector(to_signed(223,bitWidth));
      c_rom(30) <= std_logic_vector(to_signed(220,bitWidth));
      c_rom(31) <= std_logic_vector(to_signed(218,bitWidth));
      c_rom(32) <= std_logic_vector(to_signed(216,bitWidth));
      c_rom(33) <= std_logic_vector(to_signed(213,bitWidth));
      c_rom(34) <= std_logic_vector(to_signed(211,bitWidth));
      c_rom(35) <= std_logic_vector(to_signed(208,bitWidth));
      c_rom(36) <= std_logic_vector(to_signed(206,bitWidth));
      c_rom(37) <= std_logic_vector(to_signed(203,bitWidth));
      c_rom(38) <= std_logic_vector(to_signed(200,bitWidth));
      c_rom(39) <= std_logic_vector(to_signed(198,bitWidth));
      c_rom(40) <= std_logic_vector(to_signed(195,bitWidth));
      c_rom(41) <= std_logic_vector(to_signed(192,bitWidth));
      c_rom(42) <= std_logic_vector(to_signed(189,bitWidth));
      c_rom(43) <= std_logic_vector(to_signed(186,bitWidth));
      c_rom(44) <= std_logic_vector(to_signed(183,bitWidth));
      c_rom(45) <= std_logic_vector(to_signed(180,bitWidth));
      c_rom(46) <= std_logic_vector(to_signed(177,bitWidth));
      c_rom(47) <= std_logic_vector(to_signed(173,bitWidth));
      c_rom(48) <= std_logic_vector(to_signed(170,bitWidth));
      c_rom(49) <= std_logic_vector(to_signed(167,bitWidth));
      c_rom(50) <= std_logic_vector(to_signed(163,bitWidth));
      c_rom(51) <= std_logic_vector(to_signed(160,bitWidth));
      c_rom(52) <= std_logic_vector(to_signed(156,bitWidth));
      c_rom(53) <= std_logic_vector(to_signed(153,bitWidth));
      c_rom(54) <= std_logic_vector(to_signed(149,bitWidth));
      c_rom(55) <= std_logic_vector(to_signed(146,bitWidth));
      c_rom(56) <= std_logic_vector(to_signed(142,bitWidth));
      c_rom(57) <= std_logic_vector(to_signed(138,bitWidth));
      c_rom(58) <= std_logic_vector(to_signed(135,bitWidth));
      c_rom(59) <= std_logic_vector(to_signed(131,bitWidth));
      c_rom(60) <= std_logic_vector(to_signed(127,bitWidth));
      c_rom(61) <= std_logic_vector(to_signed(123,bitWidth));
      c_rom(62) <= std_logic_vector(to_signed(119,bitWidth));
      c_rom(63) <= std_logic_vector(to_signed(115,bitWidth));
      c_rom(64) <= std_logic_vector(to_signed(111,bitWidth));
      c_rom(65) <= std_logic_vector(to_signed(107,bitWidth));
      c_rom(66) <= std_logic_vector(to_signed(103,bitWidth));
      c_rom(67) <= std_logic_vector(to_signed(99,bitWidth));
      c_rom(68) <= std_logic_vector(to_signed(95,bitWidth));
      c_rom(69) <= std_logic_vector(to_signed(91,bitWidth));
      c_rom(70) <= std_logic_vector(to_signed(87,bitWidth));
      c_rom(71) <= std_logic_vector(to_signed(83,bitWidth));
      c_rom(72) <= std_logic_vector(to_signed(78,bitWidth));
      c_rom(73) <= std_logic_vector(to_signed(74,bitWidth));
      c_rom(74) <= std_logic_vector(to_signed(70,bitWidth));
      c_rom(75) <= std_logic_vector(to_signed(65,bitWidth));
      c_rom(76) <= std_logic_vector(to_signed(61,bitWidth));
      c_rom(77) <= std_logic_vector(to_signed(57,bitWidth));
      c_rom(78) <= std_logic_vector(to_signed(53,bitWidth));
      c_rom(79) <= std_logic_vector(to_signed(48,bitWidth));
      c_rom(80) <= std_logic_vector(to_signed(44,bitWidth));
      c_rom(81) <= std_logic_vector(to_signed(39,bitWidth));
      c_rom(82) <= std_logic_vector(to_signed(35,bitWidth));
      c_rom(83) <= std_logic_vector(to_signed(31,bitWidth));
      c_rom(84) <= std_logic_vector(to_signed(26,bitWidth));
      c_rom(85) <= std_logic_vector(to_signed(22,bitWidth));
      c_rom(86) <= std_logic_vector(to_signed(17,bitWidth));
      c_rom(87) <= std_logic_vector(to_signed(13,bitWidth));
      c_rom(88) <= std_logic_vector(to_signed(8,bitWidth));
      c_rom(89) <= std_logic_vector(to_signed(4,bitWidth));
      c_rom(90) <= std_logic_vector(to_signed(0,bitWidth));
      c_rom(91) <= std_logic_vector(to_signed(-4,bitWidth));
      c_rom(92) <= std_logic_vector(to_signed(-8,bitWidth));
      c_rom(93) <= std_logic_vector(to_signed(-13,bitWidth));
      c_rom(94) <= std_logic_vector(to_signed(-17,bitWidth));
      c_rom(95) <= std_logic_vector(to_signed(-22,bitWidth));
      c_rom(96) <= std_logic_vector(to_signed(-26,bitWidth));
      c_rom(97) <= std_logic_vector(to_signed(-31,bitWidth));
      c_rom(98) <= std_logic_vector(to_signed(-35,bitWidth));
      c_rom(99) <= std_logic_vector(to_signed(-39,bitWidth));
      c_rom(100) <= std_logic_vector(to_signed(-44,bitWidth));
      c_rom(101) <= std_logic_vector(to_signed(-48,bitWidth));
      c_rom(102) <= std_logic_vector(to_signed(-53,bitWidth));
      c_rom(103) <= std_logic_vector(to_signed(-57,bitWidth));
      c_rom(104) <= std_logic_vector(to_signed(-61,bitWidth));
      c_rom(105) <= std_logic_vector(to_signed(-65,bitWidth));
      c_rom(106) <= std_logic_vector(to_signed(-70,bitWidth));
      c_rom(107) <= std_logic_vector(to_signed(-74,bitWidth));
      c_rom(108) <= std_logic_vector(to_signed(-78,bitWidth));
      c_rom(109) <= std_logic_vector(to_signed(-83,bitWidth));
      c_rom(110) <= std_logic_vector(to_signed(-87,bitWidth));
      c_rom(111) <= std_logic_vector(to_signed(-91,bitWidth));
      c_rom(112) <= std_logic_vector(to_signed(-95,bitWidth));
      c_rom(113) <= std_logic_vector(to_signed(-99,bitWidth));
      c_rom(114) <= std_logic_vector(to_signed(-103,bitWidth));
      c_rom(115) <= std_logic_vector(to_signed(-107,bitWidth));
      c_rom(116) <= std_logic_vector(to_signed(-111,bitWidth));
      c_rom(117) <= std_logic_vector(to_signed(-115,bitWidth));
      c_rom(118) <= std_logic_vector(to_signed(-119,bitWidth));
      c_rom(119) <= std_logic_vector(to_signed(-123,bitWidth));
      c_rom(120) <= std_logic_vector(to_signed(-127,bitWidth));
      c_rom(121) <= std_logic_vector(to_signed(-131,bitWidth));
      c_rom(122) <= std_logic_vector(to_signed(-135,bitWidth));
      c_rom(123) <= std_logic_vector(to_signed(-138,bitWidth));
      c_rom(124) <= std_logic_vector(to_signed(-142,bitWidth));
      c_rom(125) <= std_logic_vector(to_signed(-146,bitWidth));
      c_rom(126) <= std_logic_vector(to_signed(-149,bitWidth));
      c_rom(127) <= std_logic_vector(to_signed(-153,bitWidth));
      c_rom(128) <= std_logic_vector(to_signed(-156,bitWidth));
      c_rom(129) <= std_logic_vector(to_signed(-160,bitWidth));
      c_rom(130) <= std_logic_vector(to_signed(-163,bitWidth));
      c_rom(131) <= std_logic_vector(to_signed(-167,bitWidth));
      c_rom(132) <= std_logic_vector(to_signed(-170,bitWidth));
      c_rom(133) <= std_logic_vector(to_signed(-173,bitWidth));
      c_rom(134) <= std_logic_vector(to_signed(-177,bitWidth));
      c_rom(135) <= std_logic_vector(to_signed(-180,bitWidth));
      c_rom(136) <= std_logic_vector(to_signed(-183,bitWidth));
      c_rom(137) <= std_logic_vector(to_signed(-186,bitWidth));
      c_rom(138) <= std_logic_vector(to_signed(-189,bitWidth));
      c_rom(139) <= std_logic_vector(to_signed(-192,bitWidth));
      c_rom(140) <= std_logic_vector(to_signed(-195,bitWidth));
      c_rom(141) <= std_logic_vector(to_signed(-198,bitWidth));
      c_rom(142) <= std_logic_vector(to_signed(-200,bitWidth));
      c_rom(143) <= std_logic_vector(to_signed(-203,bitWidth));
      c_rom(144) <= std_logic_vector(to_signed(-206,bitWidth));
      c_rom(145) <= std_logic_vector(to_signed(-208,bitWidth));
      c_rom(146) <= std_logic_vector(to_signed(-211,bitWidth));
      c_rom(147) <= std_logic_vector(to_signed(-213,bitWidth));
      c_rom(148) <= std_logic_vector(to_signed(-216,bitWidth));
      c_rom(149) <= std_logic_vector(to_signed(-218,bitWidth));
      c_rom(150) <= std_logic_vector(to_signed(-220,bitWidth));
      c_rom(151) <= std_logic_vector(to_signed(-223,bitWidth));
      c_rom(152) <= std_logic_vector(to_signed(-225,bitWidth));
      c_rom(153) <= std_logic_vector(to_signed(-227,bitWidth));
      c_rom(154) <= std_logic_vector(to_signed(-229,bitWidth));
      c_rom(155) <= std_logic_vector(to_signed(-231,bitWidth));
      c_rom(156) <= std_logic_vector(to_signed(-232,bitWidth));
      c_rom(157) <= std_logic_vector(to_signed(-234,bitWidth));
      c_rom(158) <= std_logic_vector(to_signed(-236,bitWidth));
      c_rom(159) <= std_logic_vector(to_signed(-238,bitWidth));
      c_rom(160) <= std_logic_vector(to_signed(-239,bitWidth));
      c_rom(161) <= std_logic_vector(to_signed(-241,bitWidth));
      c_rom(162) <= std_logic_vector(to_signed(-242,bitWidth));
      c_rom(163) <= std_logic_vector(to_signed(-243,bitWidth));
      c_rom(164) <= std_logic_vector(to_signed(-245,bitWidth));
      c_rom(165) <= std_logic_vector(to_signed(-246,bitWidth));
      c_rom(166) <= std_logic_vector(to_signed(-247,bitWidth));
      c_rom(167) <= std_logic_vector(to_signed(-248,bitWidth));
      c_rom(168) <= std_logic_vector(to_signed(-249,bitWidth));
      c_rom(169) <= std_logic_vector(to_signed(-250,bitWidth));
      c_rom(170) <= std_logic_vector(to_signed(-251,bitWidth));
      c_rom(171) <= std_logic_vector(to_signed(-251,bitWidth));
      c_rom(172) <= std_logic_vector(to_signed(-252,bitWidth));
      c_rom(173) <= std_logic_vector(to_signed(-253,bitWidth));
      c_rom(174) <= std_logic_vector(to_signed(-253,bitWidth));
      c_rom(175) <= std_logic_vector(to_signed(-254,bitWidth));
      c_rom(176) <= std_logic_vector(to_signed(-254,bitWidth));
      c_rom(177) <= std_logic_vector(to_signed(-254,bitWidth));
      c_rom(178) <= std_logic_vector(to_signed(-254,bitWidth));
      c_rom(179) <= std_logic_vector(to_signed(-254,bitWidth));
      c_rom(180) <= std_logic_vector(to_signed(-255,bitWidth));
      c_rom(181) <= std_logic_vector(to_signed(-254,bitWidth));
      c_rom(182) <= std_logic_vector(to_signed(-254,bitWidth));
      c_rom(183) <= std_logic_vector(to_signed(-254,bitWidth));
      c_rom(184) <= std_logic_vector(to_signed(-254,bitWidth));
      c_rom(185) <= std_logic_vector(to_signed(-254,bitWidth));
      c_rom(186) <= std_logic_vector(to_signed(-253,bitWidth));
      c_rom(187) <= std_logic_vector(to_signed(-253,bitWidth));
      c_rom(188) <= std_logic_vector(to_signed(-252,bitWidth));
      c_rom(189) <= std_logic_vector(to_signed(-251,bitWidth));
      c_rom(190) <= std_logic_vector(to_signed(-251,bitWidth));
      c_rom(191) <= std_logic_vector(to_signed(-250,bitWidth));
      c_rom(192) <= std_logic_vector(to_signed(-249,bitWidth));
      c_rom(193) <= std_logic_vector(to_signed(-248,bitWidth));
      c_rom(194) <= std_logic_vector(to_signed(-247,bitWidth));
      c_rom(195) <= std_logic_vector(to_signed(-246,bitWidth));
      c_rom(196) <= std_logic_vector(to_signed(-245,bitWidth));
      c_rom(197) <= std_logic_vector(to_signed(-243,bitWidth));
      c_rom(198) <= std_logic_vector(to_signed(-242,bitWidth));
      c_rom(199) <= std_logic_vector(to_signed(-241,bitWidth));
      c_rom(200) <= std_logic_vector(to_signed(-239,bitWidth));
      c_rom(201) <= std_logic_vector(to_signed(-238,bitWidth));
      c_rom(202) <= std_logic_vector(to_signed(-236,bitWidth));
      c_rom(203) <= std_logic_vector(to_signed(-234,bitWidth));
      c_rom(204) <= std_logic_vector(to_signed(-232,bitWidth));
      c_rom(205) <= std_logic_vector(to_signed(-231,bitWidth));
      c_rom(206) <= std_logic_vector(to_signed(-229,bitWidth));
      c_rom(207) <= std_logic_vector(to_signed(-227,bitWidth));
      c_rom(208) <= std_logic_vector(to_signed(-225,bitWidth));
      c_rom(209) <= std_logic_vector(to_signed(-223,bitWidth));
      c_rom(210) <= std_logic_vector(to_signed(-220,bitWidth));
      c_rom(211) <= std_logic_vector(to_signed(-218,bitWidth));
      c_rom(212) <= std_logic_vector(to_signed(-216,bitWidth));
      c_rom(213) <= std_logic_vector(to_signed(-213,bitWidth));
      c_rom(214) <= std_logic_vector(to_signed(-211,bitWidth));
      c_rom(215) <= std_logic_vector(to_signed(-208,bitWidth));
      c_rom(216) <= std_logic_vector(to_signed(-206,bitWidth));
      c_rom(217) <= std_logic_vector(to_signed(-203,bitWidth));
      c_rom(218) <= std_logic_vector(to_signed(-200,bitWidth));
      c_rom(219) <= std_logic_vector(to_signed(-198,bitWidth));
      c_rom(220) <= std_logic_vector(to_signed(-195,bitWidth));
      c_rom(221) <= std_logic_vector(to_signed(-192,bitWidth));
      c_rom(222) <= std_logic_vector(to_signed(-189,bitWidth));
      c_rom(223) <= std_logic_vector(to_signed(-186,bitWidth));
      c_rom(224) <= std_logic_vector(to_signed(-183,bitWidth));
      c_rom(225) <= std_logic_vector(to_signed(-180,bitWidth));
      c_rom(226) <= std_logic_vector(to_signed(-177,bitWidth));
      c_rom(227) <= std_logic_vector(to_signed(-173,bitWidth));
      c_rom(228) <= std_logic_vector(to_signed(-170,bitWidth));
      c_rom(229) <= std_logic_vector(to_signed(-167,bitWidth));
      c_rom(230) <= std_logic_vector(to_signed(-163,bitWidth));
      c_rom(231) <= std_logic_vector(to_signed(-160,bitWidth));
      c_rom(232) <= std_logic_vector(to_signed(-156,bitWidth));
      c_rom(233) <= std_logic_vector(to_signed(-153,bitWidth));
      c_rom(234) <= std_logic_vector(to_signed(-149,bitWidth));
      c_rom(235) <= std_logic_vector(to_signed(-146,bitWidth));
      c_rom(236) <= std_logic_vector(to_signed(-142,bitWidth));
      c_rom(237) <= std_logic_vector(to_signed(-138,bitWidth));
      c_rom(238) <= std_logic_vector(to_signed(-135,bitWidth));
      c_rom(239) <= std_logic_vector(to_signed(-131,bitWidth));
      c_rom(240) <= std_logic_vector(to_signed(-127,bitWidth));
      c_rom(241) <= std_logic_vector(to_signed(-123,bitWidth));
      c_rom(242) <= std_logic_vector(to_signed(-119,bitWidth));
      c_rom(243) <= std_logic_vector(to_signed(-115,bitWidth));
      c_rom(244) <= std_logic_vector(to_signed(-111,bitWidth));
      c_rom(245) <= std_logic_vector(to_signed(-107,bitWidth));
      c_rom(246) <= std_logic_vector(to_signed(-103,bitWidth));
      c_rom(247) <= std_logic_vector(to_signed(-99,bitWidth));
      c_rom(248) <= std_logic_vector(to_signed(-95,bitWidth));
      c_rom(249) <= std_logic_vector(to_signed(-91,bitWidth));
      c_rom(250) <= std_logic_vector(to_signed(-87,bitWidth));
      c_rom(251) <= std_logic_vector(to_signed(-83,bitWidth));
      c_rom(252) <= std_logic_vector(to_signed(-78,bitWidth));
      c_rom(253) <= std_logic_vector(to_signed(-74,bitWidth));
      c_rom(254) <= std_logic_vector(to_signed(-70,bitWidth));
      c_rom(255) <= std_logic_vector(to_signed(-65,bitWidth));
      c_rom(256) <= std_logic_vector(to_signed(-61,bitWidth));
      c_rom(257) <= std_logic_vector(to_signed(-57,bitWidth));
      c_rom(258) <= std_logic_vector(to_signed(-53,bitWidth));
      c_rom(259) <= std_logic_vector(to_signed(-48,bitWidth));
      c_rom(260) <= std_logic_vector(to_signed(-44,bitWidth));
      c_rom(261) <= std_logic_vector(to_signed(-39,bitWidth));
      c_rom(262) <= std_logic_vector(to_signed(-35,bitWidth));
      c_rom(263) <= std_logic_vector(to_signed(-31,bitWidth));
      c_rom(264) <= std_logic_vector(to_signed(-26,bitWidth));
      c_rom(265) <= std_logic_vector(to_signed(-22,bitWidth));
      c_rom(266) <= std_logic_vector(to_signed(-17,bitWidth));
      c_rom(267) <= std_logic_vector(to_signed(-13,bitWidth));
      c_rom(268) <= std_logic_vector(to_signed(-8,bitWidth));
      c_rom(269) <= std_logic_vector(to_signed(-4,bitWidth));
      c_rom(270) <= std_logic_vector(to_signed(0,bitWidth));
      c_rom(271) <= std_logic_vector(to_signed(4,bitWidth));
      c_rom(272) <= std_logic_vector(to_signed(8,bitWidth));
      c_rom(273) <= std_logic_vector(to_signed(13,bitWidth));
      c_rom(274) <= std_logic_vector(to_signed(17,bitWidth));
      c_rom(275) <= std_logic_vector(to_signed(22,bitWidth));
      c_rom(276) <= std_logic_vector(to_signed(26,bitWidth));
      c_rom(277) <= std_logic_vector(to_signed(31,bitWidth));
      c_rom(278) <= std_logic_vector(to_signed(35,bitWidth));
      c_rom(279) <= std_logic_vector(to_signed(39,bitWidth));
      c_rom(280) <= std_logic_vector(to_signed(44,bitWidth));
      c_rom(281) <= std_logic_vector(to_signed(48,bitWidth));
      c_rom(282) <= std_logic_vector(to_signed(53,bitWidth));
      c_rom(283) <= std_logic_vector(to_signed(57,bitWidth));
      c_rom(284) <= std_logic_vector(to_signed(61,bitWidth));
      c_rom(285) <= std_logic_vector(to_signed(65,bitWidth));
      c_rom(286) <= std_logic_vector(to_signed(70,bitWidth));
      c_rom(287) <= std_logic_vector(to_signed(74,bitWidth));
      c_rom(288) <= std_logic_vector(to_signed(78,bitWidth));
      c_rom(289) <= std_logic_vector(to_signed(83,bitWidth));
      c_rom(290) <= std_logic_vector(to_signed(87,bitWidth));
      c_rom(291) <= std_logic_vector(to_signed(91,bitWidth));
      c_rom(292) <= std_logic_vector(to_signed(95,bitWidth));
      c_rom(293) <= std_logic_vector(to_signed(99,bitWidth));
      c_rom(294) <= std_logic_vector(to_signed(103,bitWidth));
      c_rom(295) <= std_logic_vector(to_signed(107,bitWidth));
      c_rom(296) <= std_logic_vector(to_signed(111,bitWidth));
      c_rom(297) <= std_logic_vector(to_signed(115,bitWidth));
      c_rom(298) <= std_logic_vector(to_signed(119,bitWidth));
      c_rom(299) <= std_logic_vector(to_signed(123,bitWidth));
      c_rom(300) <= std_logic_vector(to_signed(127,bitWidth));
      c_rom(301) <= std_logic_vector(to_signed(131,bitWidth));
      c_rom(302) <= std_logic_vector(to_signed(135,bitWidth));
      c_rom(303) <= std_logic_vector(to_signed(138,bitWidth));
      c_rom(304) <= std_logic_vector(to_signed(142,bitWidth));
      c_rom(305) <= std_logic_vector(to_signed(146,bitWidth));
      c_rom(306) <= std_logic_vector(to_signed(149,bitWidth));
      c_rom(307) <= std_logic_vector(to_signed(153,bitWidth));
      c_rom(308) <= std_logic_vector(to_signed(156,bitWidth));
      c_rom(309) <= std_logic_vector(to_signed(160,bitWidth));
      c_rom(310) <= std_logic_vector(to_signed(163,bitWidth));
      c_rom(311) <= std_logic_vector(to_signed(167,bitWidth));
      c_rom(312) <= std_logic_vector(to_signed(170,bitWidth));
      c_rom(313) <= std_logic_vector(to_signed(173,bitWidth));
      c_rom(314) <= std_logic_vector(to_signed(177,bitWidth));
      c_rom(315) <= std_logic_vector(to_signed(180,bitWidth));
      c_rom(316) <= std_logic_vector(to_signed(183,bitWidth));
      c_rom(317) <= std_logic_vector(to_signed(186,bitWidth));
      c_rom(318) <= std_logic_vector(to_signed(189,bitWidth));
      c_rom(319) <= std_logic_vector(to_signed(192,bitWidth));
      c_rom(320) <= std_logic_vector(to_signed(195,bitWidth));
      c_rom(321) <= std_logic_vector(to_signed(198,bitWidth));
      c_rom(322) <= std_logic_vector(to_signed(200,bitWidth));
      c_rom(323) <= std_logic_vector(to_signed(203,bitWidth));
      c_rom(324) <= std_logic_vector(to_signed(206,bitWidth));
      c_rom(325) <= std_logic_vector(to_signed(208,bitWidth));
      c_rom(326) <= std_logic_vector(to_signed(211,bitWidth));
      c_rom(327) <= std_logic_vector(to_signed(213,bitWidth));
      c_rom(328) <= std_logic_vector(to_signed(216,bitWidth));
      c_rom(329) <= std_logic_vector(to_signed(218,bitWidth));
      c_rom(330) <= std_logic_vector(to_signed(220,bitWidth));
      c_rom(331) <= std_logic_vector(to_signed(223,bitWidth));
      c_rom(332) <= std_logic_vector(to_signed(225,bitWidth));
      c_rom(333) <= std_logic_vector(to_signed(227,bitWidth));
      c_rom(334) <= std_logic_vector(to_signed(229,bitWidth));
      c_rom(335) <= std_logic_vector(to_signed(231,bitWidth));
      c_rom(336) <= std_logic_vector(to_signed(232,bitWidth));
      c_rom(337) <= std_logic_vector(to_signed(234,bitWidth));
      c_rom(338) <= std_logic_vector(to_signed(236,bitWidth));
      c_rom(339) <= std_logic_vector(to_signed(238,bitWidth));
      c_rom(340) <= std_logic_vector(to_signed(239,bitWidth));
      c_rom(341) <= std_logic_vector(to_signed(241,bitWidth));
      c_rom(342) <= std_logic_vector(to_signed(242,bitWidth));
      c_rom(343) <= std_logic_vector(to_signed(243,bitWidth));
      c_rom(344) <= std_logic_vector(to_signed(245,bitWidth));
      c_rom(345) <= std_logic_vector(to_signed(246,bitWidth));
      c_rom(346) <= std_logic_vector(to_signed(247,bitWidth));
      c_rom(347) <= std_logic_vector(to_signed(248,bitWidth));
      c_rom(348) <= std_logic_vector(to_signed(249,bitWidth));
      c_rom(349) <= std_logic_vector(to_signed(250,bitWidth));
      c_rom(350) <= std_logic_vector(to_signed(251,bitWidth));
      c_rom(351) <= std_logic_vector(to_signed(251,bitWidth));
      c_rom(352) <= std_logic_vector(to_signed(252,bitWidth));
      c_rom(353) <= std_logic_vector(to_signed(253,bitWidth));
      c_rom(354) <= std_logic_vector(to_signed(253,bitWidth));
      c_rom(355) <= std_logic_vector(to_signed(254,bitWidth));
      c_rom(356) <= std_logic_vector(to_signed(254,bitWidth));
      c_rom(357) <= std_logic_vector(to_signed(254,bitWidth));
      c_rom(358) <= std_logic_vector(to_signed(254,bitWidth));
      c_rom(359) <= std_logic_vector(to_signed(254,bitWidth));
      c_rom(360) <= std_logic_vector(to_signed(255,bitWidth));

      end if;
    end procedure;
end package body fftpackage;