library ieee;
use ieee.std_logic_1164.all;
library work;
use work.fftpackage.all;
use ieee.numeric_std.all;

entity trigo is
    port (enable : in std_logic);
end entity;



architecture trigoo of trigo is



begin
process (enable) begin
if rising_edge(enable) then 
    sin_rom(0) <= std_logic_vector(to_signed(0,bitWidth));
    sin_rom(1) <= std_logic_vector(to_signed(4,bitWidth));
    sin_rom(2) <= std_logic_vector(to_signed(8,bitWidth));
    sin_rom(3) <= std_logic_vector(to_signed(13,bitWidth));
    sin_rom(4) <= std_logic_vector(to_signed(17,bitWidth));
    sin_rom(5) <= std_logic_vector(to_signed(22,bitWidth));
    sin_rom(6) <= std_logic_vector(to_signed(26,bitWidth));
    sin_rom(7) <= std_logic_vector(to_signed(31,bitWidth));
    sin_rom(8) <= std_logic_vector(to_signed(35,bitWidth));
    sin_rom(9) <= std_logic_vector(to_signed(39,bitWidth));
    sin_rom(10) <= std_logic_vector(to_signed(44,bitWidth));
    sin_rom(11) <= std_logic_vector(to_signed(48,bitWidth));
    sin_rom(12) <= std_logic_vector(to_signed(53,bitWidth));
    sin_rom(13) <= std_logic_vector(to_signed(57,bitWidth));
    sin_rom(14) <= std_logic_vector(to_signed(61,bitWidth));
    sin_rom(15) <= std_logic_vector(to_signed(65,bitWidth));
    sin_rom(16) <= std_logic_vector(to_signed(70,bitWidth));
    sin_rom(17) <= std_logic_vector(to_signed(74,bitWidth));
    sin_rom(18) <= std_logic_vector(to_signed(78,bitWidth));
    sin_rom(19) <= std_logic_vector(to_signed(83,bitWidth));
    sin_rom(20) <= std_logic_vector(to_signed(87,bitWidth));
    sin_rom(21) <= std_logic_vector(to_signed(91,bitWidth));
    sin_rom(22) <= std_logic_vector(to_signed(95,bitWidth));
    sin_rom(23) <= std_logic_vector(to_signed(99,bitWidth));
    sin_rom(24) <= std_logic_vector(to_signed(103,bitWidth));
    sin_rom(25) <= std_logic_vector(to_signed(107,bitWidth));
    sin_rom(26) <= std_logic_vector(to_signed(111,bitWidth));
    sin_rom(27) <= std_logic_vector(to_signed(115,bitWidth));
    sin_rom(28) <= std_logic_vector(to_signed(119,bitWidth));
    sin_rom(29) <= std_logic_vector(to_signed(123,bitWidth));
    sin_rom(30) <= std_logic_vector(to_signed(127,bitWidth));
    sin_rom(31) <= std_logic_vector(to_signed(131,bitWidth));
    sin_rom(32) <= std_logic_vector(to_signed(135,bitWidth));
    sin_rom(33) <= std_logic_vector(to_signed(138,bitWidth));
    sin_rom(34) <= std_logic_vector(to_signed(142,bitWidth));
    sin_rom(35) <= std_logic_vector(to_signed(146,bitWidth));
    sin_rom(36) <= std_logic_vector(to_signed(149,bitWidth));
    sin_rom(37) <= std_logic_vector(to_signed(153,bitWidth));
    sin_rom(38) <= std_logic_vector(to_signed(156,bitWidth));
    sin_rom(39) <= std_logic_vector(to_signed(160,bitWidth));
    sin_rom(40) <= std_logic_vector(to_signed(163,bitWidth));
    sin_rom(41) <= std_logic_vector(to_signed(167,bitWidth));
    sin_rom(42) <= std_logic_vector(to_signed(170,bitWidth));
    sin_rom(43) <= std_logic_vector(to_signed(173,bitWidth));
    sin_rom(44) <= std_logic_vector(to_signed(177,bitWidth));
    sin_rom(45) <= std_logic_vector(to_signed(180,bitWidth));
    sin_rom(46) <= std_logic_vector(to_signed(183,bitWidth));
    sin_rom(47) <= std_logic_vector(to_signed(186,bitWidth));
    sin_rom(48) <= std_logic_vector(to_signed(189,bitWidth));
    sin_rom(49) <= std_logic_vector(to_signed(192,bitWidth));
    sin_rom(50) <= std_logic_vector(to_signed(195,bitWidth));
    sin_rom(51) <= std_logic_vector(to_signed(198,bitWidth));
    sin_rom(52) <= std_logic_vector(to_signed(200,bitWidth));
    sin_rom(53) <= std_logic_vector(to_signed(203,bitWidth));
    sin_rom(54) <= std_logic_vector(to_signed(206,bitWidth));
    sin_rom(55) <= std_logic_vector(to_signed(208,bitWidth));
    sin_rom(56) <= std_logic_vector(to_signed(211,bitWidth));
    sin_rom(57) <= std_logic_vector(to_signed(213,bitWidth));
    sin_rom(58) <= std_logic_vector(to_signed(216,bitWidth));
    sin_rom(59) <= std_logic_vector(to_signed(218,bitWidth));
    sin_rom(60) <= std_logic_vector(to_signed(220,bitWidth));
    sin_rom(61) <= std_logic_vector(to_signed(223,bitWidth));
    sin_rom(62) <= std_logic_vector(to_signed(225,bitWidth));
    sin_rom(63) <= std_logic_vector(to_signed(227,bitWidth));
    sin_rom(64) <= std_logic_vector(to_signed(229,bitWidth));
    sin_rom(65) <= std_logic_vector(to_signed(231,bitWidth));
    sin_rom(66) <= std_logic_vector(to_signed(232,bitWidth));
    sin_rom(67) <= std_logic_vector(to_signed(234,bitWidth));
    sin_rom(68) <= std_logic_vector(to_signed(236,bitWidth));
    sin_rom(69) <= std_logic_vector(to_signed(238,bitWidth));
    sin_rom(70) <= std_logic_vector(to_signed(239,bitWidth));
    sin_rom(71) <= std_logic_vector(to_signed(241,bitWidth));
    sin_rom(72) <= std_logic_vector(to_signed(242,bitWidth));
    sin_rom(73) <= std_logic_vector(to_signed(243,bitWidth));
    sin_rom(74) <= std_logic_vector(to_signed(245,bitWidth));
    sin_rom(75) <= std_logic_vector(to_signed(246,bitWidth));
    sin_rom(76) <= std_logic_vector(to_signed(247,bitWidth));
    sin_rom(77) <= std_logic_vector(to_signed(248,bitWidth));
    sin_rom(78) <= std_logic_vector(to_signed(249,bitWidth));
    sin_rom(79) <= std_logic_vector(to_signed(250,bitWidth));
    sin_rom(80) <= std_logic_vector(to_signed(251,bitWidth));
    sin_rom(81) <= std_logic_vector(to_signed(251,bitWidth));
    sin_rom(82) <= std_logic_vector(to_signed(252,bitWidth));
    sin_rom(83) <= std_logic_vector(to_signed(253,bitWidth));
    sin_rom(84) <= std_logic_vector(to_signed(253,bitWidth));
    sin_rom(85) <= std_logic_vector(to_signed(254,bitWidth));
    sin_rom(86) <= std_logic_vector(to_signed(254,bitWidth));
    sin_rom(87) <= std_logic_vector(to_signed(254,bitWidth));
    sin_rom(88) <= std_logic_vector(to_signed(254,bitWidth));
    sin_rom(89) <= std_logic_vector(to_signed(254,bitWidth));
    sin_rom(90) <= std_logic_vector(to_signed(255,bitWidth));
    sin_rom(91) <= std_logic_vector(to_signed(254,bitWidth));
    sin_rom(92) <= std_logic_vector(to_signed(254,bitWidth));
    sin_rom(93) <= std_logic_vector(to_signed(254,bitWidth));
    sin_rom(94) <= std_logic_vector(to_signed(254,bitWidth));
    sin_rom(95) <= std_logic_vector(to_signed(254,bitWidth));
    sin_rom(96) <= std_logic_vector(to_signed(253,bitWidth));
    sin_rom(97) <= std_logic_vector(to_signed(253,bitWidth));
    sin_rom(98) <= std_logic_vector(to_signed(252,bitWidth));
    sin_rom(99) <= std_logic_vector(to_signed(251,bitWidth));
    sin_rom(100) <= std_logic_vector(to_signed(251,bitWidth));
    sin_rom(101) <= std_logic_vector(to_signed(250,bitWidth));
    sin_rom(102) <= std_logic_vector(to_signed(249,bitWidth));
    sin_rom(103) <= std_logic_vector(to_signed(248,bitWidth));
    sin_rom(104) <= std_logic_vector(to_signed(247,bitWidth));
    sin_rom(105) <= std_logic_vector(to_signed(246,bitWidth));
    sin_rom(106) <= std_logic_vector(to_signed(245,bitWidth));
    sin_rom(107) <= std_logic_vector(to_signed(243,bitWidth));
    sin_rom(108) <= std_logic_vector(to_signed(242,bitWidth));
    sin_rom(109) <= std_logic_vector(to_signed(241,bitWidth));
    sin_rom(110) <= std_logic_vector(to_signed(239,bitWidth));
    sin_rom(111) <= std_logic_vector(to_signed(238,bitWidth));
    sin_rom(112) <= std_logic_vector(to_signed(236,bitWidth));
    sin_rom(113) <= std_logic_vector(to_signed(234,bitWidth));
    sin_rom(114) <= std_logic_vector(to_signed(232,bitWidth));
    sin_rom(115) <= std_logic_vector(to_signed(231,bitWidth));
    sin_rom(116) <= std_logic_vector(to_signed(229,bitWidth));
    sin_rom(117) <= std_logic_vector(to_signed(227,bitWidth));
    sin_rom(118) <= std_logic_vector(to_signed(225,bitWidth));
    sin_rom(119) <= std_logic_vector(to_signed(223,bitWidth));
    sin_rom(120) <= std_logic_vector(to_signed(220,bitWidth));
    sin_rom(121) <= std_logic_vector(to_signed(218,bitWidth));
    sin_rom(122) <= std_logic_vector(to_signed(216,bitWidth));
    sin_rom(123) <= std_logic_vector(to_signed(213,bitWidth));
    sin_rom(124) <= std_logic_vector(to_signed(211,bitWidth));
    sin_rom(125) <= std_logic_vector(to_signed(208,bitWidth));
    sin_rom(126) <= std_logic_vector(to_signed(206,bitWidth));
    sin_rom(127) <= std_logic_vector(to_signed(203,bitWidth));
    sin_rom(128) <= std_logic_vector(to_signed(200,bitWidth));
    sin_rom(129) <= std_logic_vector(to_signed(198,bitWidth));
    sin_rom(130) <= std_logic_vector(to_signed(195,bitWidth));
    sin_rom(131) <= std_logic_vector(to_signed(192,bitWidth));
    sin_rom(132) <= std_logic_vector(to_signed(189,bitWidth));
    sin_rom(133) <= std_logic_vector(to_signed(186,bitWidth));
    sin_rom(134) <= std_logic_vector(to_signed(183,bitWidth));
    sin_rom(135) <= std_logic_vector(to_signed(180,bitWidth));
    sin_rom(136) <= std_logic_vector(to_signed(177,bitWidth));
    sin_rom(137) <= std_logic_vector(to_signed(173,bitWidth));
    sin_rom(138) <= std_logic_vector(to_signed(170,bitWidth));
    sin_rom(139) <= std_logic_vector(to_signed(167,bitWidth));
    sin_rom(140) <= std_logic_vector(to_signed(163,bitWidth));
    sin_rom(141) <= std_logic_vector(to_signed(160,bitWidth));
    sin_rom(142) <= std_logic_vector(to_signed(156,bitWidth));
    sin_rom(143) <= std_logic_vector(to_signed(153,bitWidth));
    sin_rom(144) <= std_logic_vector(to_signed(149,bitWidth));
    sin_rom(145) <= std_logic_vector(to_signed(146,bitWidth));
    sin_rom(146) <= std_logic_vector(to_signed(142,bitWidth));
    sin_rom(147) <= std_logic_vector(to_signed(138,bitWidth));
    sin_rom(148) <= std_logic_vector(to_signed(135,bitWidth));
    sin_rom(149) <= std_logic_vector(to_signed(131,bitWidth));
    sin_rom(150) <= std_logic_vector(to_signed(127,bitWidth));
    sin_rom(151) <= std_logic_vector(to_signed(123,bitWidth));
    sin_rom(152) <= std_logic_vector(to_signed(119,bitWidth));
    sin_rom(153) <= std_logic_vector(to_signed(115,bitWidth));
    sin_rom(154) <= std_logic_vector(to_signed(111,bitWidth));
    sin_rom(155) <= std_logic_vector(to_signed(107,bitWidth));
    sin_rom(156) <= std_logic_vector(to_signed(103,bitWidth));
    sin_rom(157) <= std_logic_vector(to_signed(99,bitWidth));
    sin_rom(158) <= std_logic_vector(to_signed(95,bitWidth));
    sin_rom(159) <= std_logic_vector(to_signed(91,bitWidth));
    sin_rom(160) <= std_logic_vector(to_signed(87,bitWidth));
    sin_rom(161) <= std_logic_vector(to_signed(83,bitWidth));
    sin_rom(162) <= std_logic_vector(to_signed(78,bitWidth));
    sin_rom(163) <= std_logic_vector(to_signed(74,bitWidth));
    sin_rom(164) <= std_logic_vector(to_signed(70,bitWidth));
    sin_rom(165) <= std_logic_vector(to_signed(65,bitWidth));
    sin_rom(166) <= std_logic_vector(to_signed(61,bitWidth));
    sin_rom(167) <= std_logic_vector(to_signed(57,bitWidth));
    sin_rom(168) <= std_logic_vector(to_signed(53,bitWidth));
    sin_rom(169) <= std_logic_vector(to_signed(48,bitWidth));
    sin_rom(170) <= std_logic_vector(to_signed(44,bitWidth));
    sin_rom(171) <= std_logic_vector(to_signed(39,bitWidth));
    sin_rom(172) <= std_logic_vector(to_signed(35,bitWidth));
    sin_rom(173) <= std_logic_vector(to_signed(31,bitWidth));
    sin_rom(174) <= std_logic_vector(to_signed(26,bitWidth));
    sin_rom(175) <= std_logic_vector(to_signed(22,bitWidth));
    sin_rom(176) <= std_logic_vector(to_signed(17,bitWidth));
    sin_rom(177) <= std_logic_vector(to_signed(13,bitWidth));
    sin_rom(178) <= std_logic_vector(to_signed(8,bitWidth));
    sin_rom(179) <= std_logic_vector(to_signed(4,bitWidth));
    sin_rom(180) <= std_logic_vector(to_signed(0,bitWidth));
    sin_rom(181) <= std_logic_vector(to_signed(-4,bitWidth));
    sin_rom(182) <= std_logic_vector(to_signed(-8,bitWidth));
    sin_rom(183) <= std_logic_vector(to_signed(-13,bitWidth));
    sin_rom(184) <= std_logic_vector(to_signed(-17,bitWidth));
    sin_rom(185) <= std_logic_vector(to_signed(-22,bitWidth));
    sin_rom(186) <= std_logic_vector(to_signed(-26,bitWidth));
    sin_rom(187) <= std_logic_vector(to_signed(-31,bitWidth));
    sin_rom(188) <= std_logic_vector(to_signed(-35,bitWidth));
    sin_rom(189) <= std_logic_vector(to_signed(-39,bitWidth));
    sin_rom(190) <= std_logic_vector(to_signed(-44,bitWidth));
    sin_rom(191) <= std_logic_vector(to_signed(-48,bitWidth));
    sin_rom(192) <= std_logic_vector(to_signed(-53,bitWidth));
    sin_rom(193) <= std_logic_vector(to_signed(-57,bitWidth));
    sin_rom(194) <= std_logic_vector(to_signed(-61,bitWidth));
    sin_rom(195) <= std_logic_vector(to_signed(-65,bitWidth));
    sin_rom(196) <= std_logic_vector(to_signed(-70,bitWidth));
    sin_rom(197) <= std_logic_vector(to_signed(-74,bitWidth));
    sin_rom(198) <= std_logic_vector(to_signed(-78,bitWidth));
    sin_rom(199) <= std_logic_vector(to_signed(-83,bitWidth));
    sin_rom(200) <= std_logic_vector(to_signed(-87,bitWidth));
    sin_rom(201) <= std_logic_vector(to_signed(-91,bitWidth));
    sin_rom(202) <= std_logic_vector(to_signed(-95,bitWidth));
    sin_rom(203) <= std_logic_vector(to_signed(-99,bitWidth));
    sin_rom(204) <= std_logic_vector(to_signed(-103,bitWidth));
    sin_rom(205) <= std_logic_vector(to_signed(-107,bitWidth));
    sin_rom(206) <= std_logic_vector(to_signed(-111,bitWidth));
    sin_rom(207) <= std_logic_vector(to_signed(-115,bitWidth));
    sin_rom(208) <= std_logic_vector(to_signed(-119,bitWidth));
    sin_rom(209) <= std_logic_vector(to_signed(-123,bitWidth));
    sin_rom(210) <= std_logic_vector(to_signed(-127,bitWidth));
    sin_rom(211) <= std_logic_vector(to_signed(-131,bitWidth));
    sin_rom(212) <= std_logic_vector(to_signed(-135,bitWidth));
    sin_rom(213) <= std_logic_vector(to_signed(-138,bitWidth));
    sin_rom(214) <= std_logic_vector(to_signed(-142,bitWidth));
    sin_rom(215) <= std_logic_vector(to_signed(-146,bitWidth));
    sin_rom(216) <= std_logic_vector(to_signed(-149,bitWidth));
    sin_rom(217) <= std_logic_vector(to_signed(-153,bitWidth));
    sin_rom(218) <= std_logic_vector(to_signed(-156,bitWidth));
    sin_rom(219) <= std_logic_vector(to_signed(-160,bitWidth));
    sin_rom(220) <= std_logic_vector(to_signed(-163,bitWidth));
    sin_rom(221) <= std_logic_vector(to_signed(-167,bitWidth));
    sin_rom(222) <= std_logic_vector(to_signed(-170,bitWidth));
    sin_rom(223) <= std_logic_vector(to_signed(-173,bitWidth));
    sin_rom(224) <= std_logic_vector(to_signed(-177,bitWidth));
    sin_rom(225) <= std_logic_vector(to_signed(-180,bitWidth));
    sin_rom(226) <= std_logic_vector(to_signed(-183,bitWidth));
    sin_rom(227) <= std_logic_vector(to_signed(-186,bitWidth));
    sin_rom(228) <= std_logic_vector(to_signed(-189,bitWidth));
    sin_rom(229) <= std_logic_vector(to_signed(-192,bitWidth));
    sin_rom(230) <= std_logic_vector(to_signed(-195,bitWidth));
    sin_rom(231) <= std_logic_vector(to_signed(-198,bitWidth));
    sin_rom(232) <= std_logic_vector(to_signed(-200,bitWidth));
    sin_rom(233) <= std_logic_vector(to_signed(-203,bitWidth));
    sin_rom(234) <= std_logic_vector(to_signed(-206,bitWidth));
    sin_rom(235) <= std_logic_vector(to_signed(-208,bitWidth));
    sin_rom(236) <= std_logic_vector(to_signed(-211,bitWidth));
    sin_rom(237) <= std_logic_vector(to_signed(-213,bitWidth));
    sin_rom(238) <= std_logic_vector(to_signed(-216,bitWidth));
    sin_rom(239) <= std_logic_vector(to_signed(-218,bitWidth));
    sin_rom(240) <= std_logic_vector(to_signed(-220,bitWidth));
    sin_rom(241) <= std_logic_vector(to_signed(-223,bitWidth));
    sin_rom(242) <= std_logic_vector(to_signed(-225,bitWidth));
    sin_rom(243) <= std_logic_vector(to_signed(-227,bitWidth));
    sin_rom(244) <= std_logic_vector(to_signed(-229,bitWidth));
    sin_rom(245) <= std_logic_vector(to_signed(-231,bitWidth));
    sin_rom(246) <= std_logic_vector(to_signed(-232,bitWidth));
    sin_rom(247) <= std_logic_vector(to_signed(-234,bitWidth));
    sin_rom(248) <= std_logic_vector(to_signed(-236,bitWidth));
    sin_rom(249) <= std_logic_vector(to_signed(-238,bitWidth));
    sin_rom(250) <= std_logic_vector(to_signed(-239,bitWidth));
    sin_rom(251) <= std_logic_vector(to_signed(-241,bitWidth));
    sin_rom(252) <= std_logic_vector(to_signed(-242,bitWidth));
    sin_rom(253) <= std_logic_vector(to_signed(-243,bitWidth));
    sin_rom(254) <= std_logic_vector(to_signed(-245,bitWidth));
    sin_rom(255) <= std_logic_vector(to_signed(-246,bitWidth));
    sin_rom(256) <= std_logic_vector(to_signed(-247,bitWidth));
    sin_rom(257) <= std_logic_vector(to_signed(-248,bitWidth));
    sin_rom(258) <= std_logic_vector(to_signed(-249,bitWidth));
    sin_rom(259) <= std_logic_vector(to_signed(-250,bitWidth));
    sin_rom(260) <= std_logic_vector(to_signed(-251,bitWidth));
    sin_rom(261) <= std_logic_vector(to_signed(-251,bitWidth));
    sin_rom(262) <= std_logic_vector(to_signed(-252,bitWidth));
    sin_rom(263) <= std_logic_vector(to_signed(-253,bitWidth));
    sin_rom(264) <= std_logic_vector(to_signed(-253,bitWidth));
    sin_rom(265) <= std_logic_vector(to_signed(-254,bitWidth));
    sin_rom(266) <= std_logic_vector(to_signed(-254,bitWidth));
    sin_rom(267) <= std_logic_vector(to_signed(-254,bitWidth));
    sin_rom(268) <= std_logic_vector(to_signed(-254,bitWidth));
    sin_rom(269) <= std_logic_vector(to_signed(-254,bitWidth));
    sin_rom(270) <= std_logic_vector(to_signed(-255,bitWidth));
    sin_rom(271) <= std_logic_vector(to_signed(-254,bitWidth));
    sin_rom(272) <= std_logic_vector(to_signed(-254,bitWidth));
    sin_rom(273) <= std_logic_vector(to_signed(-254,bitWidth));
    sin_rom(274) <= std_logic_vector(to_signed(-254,bitWidth));
    sin_rom(275) <= std_logic_vector(to_signed(-254,bitWidth));
    sin_rom(276) <= std_logic_vector(to_signed(-253,bitWidth));
    sin_rom(277) <= std_logic_vector(to_signed(-253,bitWidth));
    sin_rom(278) <= std_logic_vector(to_signed(-252,bitWidth));
    sin_rom(279) <= std_logic_vector(to_signed(-251,bitWidth));
    sin_rom(280) <= std_logic_vector(to_signed(-251,bitWidth));
    sin_rom(281) <= std_logic_vector(to_signed(-250,bitWidth));
    sin_rom(282) <= std_logic_vector(to_signed(-249,bitWidth));
    sin_rom(283) <= std_logic_vector(to_signed(-248,bitWidth));
    sin_rom(284) <= std_logic_vector(to_signed(-247,bitWidth));
    sin_rom(285) <= std_logic_vector(to_signed(-246,bitWidth));
    sin_rom(286) <= std_logic_vector(to_signed(-245,bitWidth));
    sin_rom(287) <= std_logic_vector(to_signed(-243,bitWidth));
    sin_rom(288) <= std_logic_vector(to_signed(-242,bitWidth));
    sin_rom(289) <= std_logic_vector(to_signed(-241,bitWidth));
    sin_rom(290) <= std_logic_vector(to_signed(-239,bitWidth));
    sin_rom(291) <= std_logic_vector(to_signed(-238,bitWidth));
    sin_rom(292) <= std_logic_vector(to_signed(-236,bitWidth));
    sin_rom(293) <= std_logic_vector(to_signed(-234,bitWidth));
    sin_rom(294) <= std_logic_vector(to_signed(-232,bitWidth));
    sin_rom(295) <= std_logic_vector(to_signed(-231,bitWidth));
    sin_rom(296) <= std_logic_vector(to_signed(-229,bitWidth));
    sin_rom(297) <= std_logic_vector(to_signed(-227,bitWidth));
    sin_rom(298) <= std_logic_vector(to_signed(-225,bitWidth));
    sin_rom(299) <= std_logic_vector(to_signed(-223,bitWidth));
    sin_rom(300) <= std_logic_vector(to_signed(-220,bitWidth));
    sin_rom(301) <= std_logic_vector(to_signed(-218,bitWidth));
    sin_rom(302) <= std_logic_vector(to_signed(-216,bitWidth));
    sin_rom(303) <= std_logic_vector(to_signed(-213,bitWidth));
    sin_rom(304) <= std_logic_vector(to_signed(-211,bitWidth));
    sin_rom(305) <= std_logic_vector(to_signed(-208,bitWidth));
    sin_rom(306) <= std_logic_vector(to_signed(-206,bitWidth));
    sin_rom(307) <= std_logic_vector(to_signed(-203,bitWidth));
    sin_rom(308) <= std_logic_vector(to_signed(-200,bitWidth));
    sin_rom(309) <= std_logic_vector(to_signed(-198,bitWidth));
    sin_rom(310) <= std_logic_vector(to_signed(-195,bitWidth));
    sin_rom(311) <= std_logic_vector(to_signed(-192,bitWidth));
    sin_rom(312) <= std_logic_vector(to_signed(-189,bitWidth));
    sin_rom(313) <= std_logic_vector(to_signed(-186,bitWidth));
    sin_rom(314) <= std_logic_vector(to_signed(-183,bitWidth));
    sin_rom(315) <= std_logic_vector(to_signed(-180,bitWidth));
    sin_rom(316) <= std_logic_vector(to_signed(-177,bitWidth));
    sin_rom(317) <= std_logic_vector(to_signed(-173,bitWidth));
    sin_rom(318) <= std_logic_vector(to_signed(-170,bitWidth));
    sin_rom(319) <= std_logic_vector(to_signed(-167,bitWidth));
    sin_rom(320) <= std_logic_vector(to_signed(-163,bitWidth));
    sin_rom(321) <= std_logic_vector(to_signed(-160,bitWidth));
    sin_rom(322) <= std_logic_vector(to_signed(-156,bitWidth));
    sin_rom(323) <= std_logic_vector(to_signed(-153,bitWidth));
    sin_rom(324) <= std_logic_vector(to_signed(-149,bitWidth));
    sin_rom(325) <= std_logic_vector(to_signed(-146,bitWidth));
    sin_rom(326) <= std_logic_vector(to_signed(-142,bitWidth));
    sin_rom(327) <= std_logic_vector(to_signed(-138,bitWidth));
    sin_rom(328) <= std_logic_vector(to_signed(-135,bitWidth));
    sin_rom(329) <= std_logic_vector(to_signed(-131,bitWidth));
    sin_rom(330) <= std_logic_vector(to_signed(-127,bitWidth));
    sin_rom(331) <= std_logic_vector(to_signed(-123,bitWidth));
    sin_rom(332) <= std_logic_vector(to_signed(-119,bitWidth));
    sin_rom(333) <= std_logic_vector(to_signed(-115,bitWidth));
    sin_rom(334) <= std_logic_vector(to_signed(-111,bitWidth));
    sin_rom(335) <= std_logic_vector(to_signed(-107,bitWidth));
    sin_rom(336) <= std_logic_vector(to_signed(-103,bitWidth));
    sin_rom(337) <= std_logic_vector(to_signed(-99,bitWidth));
    sin_rom(338) <= std_logic_vector(to_signed(-95,bitWidth));
    sin_rom(339) <= std_logic_vector(to_signed(-91,bitWidth));
    sin_rom(340) <= std_logic_vector(to_signed(-87,bitWidth));
    sin_rom(341) <= std_logic_vector(to_signed(-83,bitWidth));
    sin_rom(342) <= std_logic_vector(to_signed(-78,bitWidth));
    sin_rom(343) <= std_logic_vector(to_signed(-74,bitWidth));
    sin_rom(344) <= std_logic_vector(to_signed(-70,bitWidth));
    sin_rom(345) <= std_logic_vector(to_signed(-65,bitWidth));
    sin_rom(346) <= std_logic_vector(to_signed(-61,bitWidth));
    sin_rom(347) <= std_logic_vector(to_signed(-57,bitWidth));
    sin_rom(348) <= std_logic_vector(to_signed(-53,bitWidth));
    sin_rom(349) <= std_logic_vector(to_signed(-48,bitWidth));
    sin_rom(350) <= std_logic_vector(to_signed(-44,bitWidth));
    sin_rom(351) <= std_logic_vector(to_signed(-39,bitWidth));
    sin_rom(352) <= std_logic_vector(to_signed(-35,bitWidth));
    sin_rom(353) <= std_logic_vector(to_signed(-31,bitWidth));
    sin_rom(354) <= std_logic_vector(to_signed(-26,bitWidth));
    sin_rom(355) <= std_logic_vector(to_signed(-22,bitWidth));
    sin_rom(356) <= std_logic_vector(to_signed(-17,bitWidth));
    sin_rom(357) <= std_logic_vector(to_signed(-13,bitWidth));
    sin_rom(358) <= std_logic_vector(to_signed(-8,bitWidth));
    sin_rom(359) <= std_logic_vector(to_signed(-4,bitWidth));
    sin_rom(360) <= std_logic_vector(to_signed(0,bitWidth));

    cos_rom(0) <= std_logic_vector(to_signed(255,bitWidth));
    cos_rom(1) <= std_logic_vector(to_signed(254,bitWidth));
    cos_rom(2) <= std_logic_vector(to_signed(254,bitWidth));
    cos_rom(3) <= std_logic_vector(to_signed(254,bitWidth));
    cos_rom(4) <= std_logic_vector(to_signed(254,bitWidth));
    cos_rom(5) <= std_logic_vector(to_signed(254,bitWidth));
    cos_rom(6) <= std_logic_vector(to_signed(253,bitWidth));
    cos_rom(7) <= std_logic_vector(to_signed(253,bitWidth));
    cos_rom(8) <= std_logic_vector(to_signed(252,bitWidth));
    cos_rom(9) <= std_logic_vector(to_signed(251,bitWidth));
    cos_rom(10) <= std_logic_vector(to_signed(251,bitWidth));
    cos_rom(11) <= std_logic_vector(to_signed(250,bitWidth));
    cos_rom(12) <= std_logic_vector(to_signed(249,bitWidth));
    cos_rom(13) <= std_logic_vector(to_signed(248,bitWidth));
    cos_rom(14) <= std_logic_vector(to_signed(247,bitWidth));
    cos_rom(15) <= std_logic_vector(to_signed(246,bitWidth));
    cos_rom(16) <= std_logic_vector(to_signed(245,bitWidth));
    cos_rom(17) <= std_logic_vector(to_signed(243,bitWidth));
    cos_rom(18) <= std_logic_vector(to_signed(242,bitWidth));
    cos_rom(19) <= std_logic_vector(to_signed(241,bitWidth));
    cos_rom(20) <= std_logic_vector(to_signed(239,bitWidth));
    cos_rom(21) <= std_logic_vector(to_signed(238,bitWidth));
    cos_rom(22) <= std_logic_vector(to_signed(236,bitWidth));
    cos_rom(23) <= std_logic_vector(to_signed(234,bitWidth));
    cos_rom(24) <= std_logic_vector(to_signed(232,bitWidth));
    cos_rom(25) <= std_logic_vector(to_signed(231,bitWidth));
    cos_rom(26) <= std_logic_vector(to_signed(229,bitWidth));
    cos_rom(27) <= std_logic_vector(to_signed(227,bitWidth));
    cos_rom(28) <= std_logic_vector(to_signed(225,bitWidth));
    cos_rom(29) <= std_logic_vector(to_signed(223,bitWidth));
    cos_rom(30) <= std_logic_vector(to_signed(220,bitWidth));
    cos_rom(31) <= std_logic_vector(to_signed(218,bitWidth));
    cos_rom(32) <= std_logic_vector(to_signed(216,bitWidth));
    cos_rom(33) <= std_logic_vector(to_signed(213,bitWidth));
    cos_rom(34) <= std_logic_vector(to_signed(211,bitWidth));
    cos_rom(35) <= std_logic_vector(to_signed(208,bitWidth));
    cos_rom(36) <= std_logic_vector(to_signed(206,bitWidth));
    cos_rom(37) <= std_logic_vector(to_signed(203,bitWidth));
    cos_rom(38) <= std_logic_vector(to_signed(200,bitWidth));
    cos_rom(39) <= std_logic_vector(to_signed(198,bitWidth));
    cos_rom(40) <= std_logic_vector(to_signed(195,bitWidth));
    cos_rom(41) <= std_logic_vector(to_signed(192,bitWidth));
    cos_rom(42) <= std_logic_vector(to_signed(189,bitWidth));
    cos_rom(43) <= std_logic_vector(to_signed(186,bitWidth));
    cos_rom(44) <= std_logic_vector(to_signed(183,bitWidth));
    cos_rom(45) <= std_logic_vector(to_signed(180,bitWidth));
    cos_rom(46) <= std_logic_vector(to_signed(177,bitWidth));
    cos_rom(47) <= std_logic_vector(to_signed(173,bitWidth));
    cos_rom(48) <= std_logic_vector(to_signed(170,bitWidth));
    cos_rom(49) <= std_logic_vector(to_signed(167,bitWidth));
    cos_rom(50) <= std_logic_vector(to_signed(163,bitWidth));
    cos_rom(51) <= std_logic_vector(to_signed(160,bitWidth));
    cos_rom(52) <= std_logic_vector(to_signed(156,bitWidth));
    cos_rom(53) <= std_logic_vector(to_signed(153,bitWidth));
    cos_rom(54) <= std_logic_vector(to_signed(149,bitWidth));
    cos_rom(55) <= std_logic_vector(to_signed(146,bitWidth));
    cos_rom(56) <= std_logic_vector(to_signed(142,bitWidth));
    cos_rom(57) <= std_logic_vector(to_signed(138,bitWidth));
    cos_rom(58) <= std_logic_vector(to_signed(135,bitWidth));
    cos_rom(59) <= std_logic_vector(to_signed(131,bitWidth));
    cos_rom(60) <= std_logic_vector(to_signed(127,bitWidth));
    cos_rom(61) <= std_logic_vector(to_signed(123,bitWidth));
    cos_rom(62) <= std_logic_vector(to_signed(119,bitWidth));
    cos_rom(63) <= std_logic_vector(to_signed(115,bitWidth));
    cos_rom(64) <= std_logic_vector(to_signed(111,bitWidth));
    cos_rom(65) <= std_logic_vector(to_signed(107,bitWidth));
    cos_rom(66) <= std_logic_vector(to_signed(103,bitWidth));
    cos_rom(67) <= std_logic_vector(to_signed(99,bitWidth));
    cos_rom(68) <= std_logic_vector(to_signed(95,bitWidth));
    cos_rom(69) <= std_logic_vector(to_signed(91,bitWidth));
    cos_rom(70) <= std_logic_vector(to_signed(87,bitWidth));
    cos_rom(71) <= std_logic_vector(to_signed(83,bitWidth));
    cos_rom(72) <= std_logic_vector(to_signed(78,bitWidth));
    cos_rom(73) <= std_logic_vector(to_signed(74,bitWidth));
    cos_rom(74) <= std_logic_vector(to_signed(70,bitWidth));
    cos_rom(75) <= std_logic_vector(to_signed(65,bitWidth));
    cos_rom(76) <= std_logic_vector(to_signed(61,bitWidth));
    cos_rom(77) <= std_logic_vector(to_signed(57,bitWidth));
    cos_rom(78) <= std_logic_vector(to_signed(53,bitWidth));
    cos_rom(79) <= std_logic_vector(to_signed(48,bitWidth));
    cos_rom(80) <= std_logic_vector(to_signed(44,bitWidth));
    cos_rom(81) <= std_logic_vector(to_signed(39,bitWidth));
    cos_rom(82) <= std_logic_vector(to_signed(35,bitWidth));
    cos_rom(83) <= std_logic_vector(to_signed(31,bitWidth));
    cos_rom(84) <= std_logic_vector(to_signed(26,bitWidth));
    cos_rom(85) <= std_logic_vector(to_signed(22,bitWidth));
    cos_rom(86) <= std_logic_vector(to_signed(17,bitWidth));
    cos_rom(87) <= std_logic_vector(to_signed(13,bitWidth));
    cos_rom(88) <= std_logic_vector(to_signed(8,bitWidth));
    cos_rom(89) <= std_logic_vector(to_signed(4,bitWidth));
    cos_rom(90) <= std_logic_vector(to_signed(0,bitWidth));
    cos_rom(91) <= std_logic_vector(to_signed(-4,bitWidth));
    cos_rom(92) <= std_logic_vector(to_signed(-8,bitWidth));
    cos_rom(93) <= std_logic_vector(to_signed(-13,bitWidth));
    cos_rom(94) <= std_logic_vector(to_signed(-17,bitWidth));
    cos_rom(95) <= std_logic_vector(to_signed(-22,bitWidth));
    cos_rom(96) <= std_logic_vector(to_signed(-26,bitWidth));
    cos_rom(97) <= std_logic_vector(to_signed(-31,bitWidth));
    cos_rom(98) <= std_logic_vector(to_signed(-35,bitWidth));
    cos_rom(99) <= std_logic_vector(to_signed(-39,bitWidth));
    cos_rom(100) <= std_logic_vector(to_signed(-44,bitWidth));
    cos_rom(101) <= std_logic_vector(to_signed(-48,bitWidth));
    cos_rom(102) <= std_logic_vector(to_signed(-53,bitWidth));
    cos_rom(103) <= std_logic_vector(to_signed(-57,bitWidth));
    cos_rom(104) <= std_logic_vector(to_signed(-61,bitWidth));
    cos_rom(105) <= std_logic_vector(to_signed(-65,bitWidth));
    cos_rom(106) <= std_logic_vector(to_signed(-70,bitWidth));
    cos_rom(107) <= std_logic_vector(to_signed(-74,bitWidth));
    cos_rom(108) <= std_logic_vector(to_signed(-78,bitWidth));
    cos_rom(109) <= std_logic_vector(to_signed(-83,bitWidth));
    cos_rom(110) <= std_logic_vector(to_signed(-87,bitWidth));
    cos_rom(111) <= std_logic_vector(to_signed(-91,bitWidth));
    cos_rom(112) <= std_logic_vector(to_signed(-95,bitWidth));
    cos_rom(113) <= std_logic_vector(to_signed(-99,bitWidth));
    cos_rom(114) <= std_logic_vector(to_signed(-103,bitWidth));
    cos_rom(115) <= std_logic_vector(to_signed(-107,bitWidth));
    cos_rom(116) <= std_logic_vector(to_signed(-111,bitWidth));
    cos_rom(117) <= std_logic_vector(to_signed(-115,bitWidth));
    cos_rom(118) <= std_logic_vector(to_signed(-119,bitWidth));
    cos_rom(119) <= std_logic_vector(to_signed(-123,bitWidth));
    cos_rom(120) <= std_logic_vector(to_signed(-127,bitWidth));
    cos_rom(121) <= std_logic_vector(to_signed(-131,bitWidth));
    cos_rom(122) <= std_logic_vector(to_signed(-135,bitWidth));
    cos_rom(123) <= std_logic_vector(to_signed(-138,bitWidth));
    cos_rom(124) <= std_logic_vector(to_signed(-142,bitWidth));
    cos_rom(125) <= std_logic_vector(to_signed(-146,bitWidth));
    cos_rom(126) <= std_logic_vector(to_signed(-149,bitWidth));
    cos_rom(127) <= std_logic_vector(to_signed(-153,bitWidth));
    cos_rom(128) <= std_logic_vector(to_signed(-156,bitWidth));
    cos_rom(129) <= std_logic_vector(to_signed(-160,bitWidth));
    cos_rom(130) <= std_logic_vector(to_signed(-163,bitWidth));
    cos_rom(131) <= std_logic_vector(to_signed(-167,bitWidth));
    cos_rom(132) <= std_logic_vector(to_signed(-170,bitWidth));
    cos_rom(133) <= std_logic_vector(to_signed(-173,bitWidth));
    cos_rom(134) <= std_logic_vector(to_signed(-177,bitWidth));
    cos_rom(135) <= std_logic_vector(to_signed(-180,bitWidth));
    cos_rom(136) <= std_logic_vector(to_signed(-183,bitWidth));
    cos_rom(137) <= std_logic_vector(to_signed(-186,bitWidth));
    cos_rom(138) <= std_logic_vector(to_signed(-189,bitWidth));
    cos_rom(139) <= std_logic_vector(to_signed(-192,bitWidth));
    cos_rom(140) <= std_logic_vector(to_signed(-195,bitWidth));
    cos_rom(141) <= std_logic_vector(to_signed(-198,bitWidth));
    cos_rom(142) <= std_logic_vector(to_signed(-200,bitWidth));
    cos_rom(143) <= std_logic_vector(to_signed(-203,bitWidth));
    cos_rom(144) <= std_logic_vector(to_signed(-206,bitWidth));
    cos_rom(145) <= std_logic_vector(to_signed(-208,bitWidth));
    cos_rom(146) <= std_logic_vector(to_signed(-211,bitWidth));
    cos_rom(147) <= std_logic_vector(to_signed(-213,bitWidth));
    cos_rom(148) <= std_logic_vector(to_signed(-216,bitWidth));
    cos_rom(149) <= std_logic_vector(to_signed(-218,bitWidth));
    cos_rom(150) <= std_logic_vector(to_signed(-220,bitWidth));
    cos_rom(151) <= std_logic_vector(to_signed(-223,bitWidth));
    cos_rom(152) <= std_logic_vector(to_signed(-225,bitWidth));
    cos_rom(153) <= std_logic_vector(to_signed(-227,bitWidth));
    cos_rom(154) <= std_logic_vector(to_signed(-229,bitWidth));
    cos_rom(155) <= std_logic_vector(to_signed(-231,bitWidth));
    cos_rom(156) <= std_logic_vector(to_signed(-232,bitWidth));
    cos_rom(157) <= std_logic_vector(to_signed(-234,bitWidth));
    cos_rom(158) <= std_logic_vector(to_signed(-236,bitWidth));
    cos_rom(159) <= std_logic_vector(to_signed(-238,bitWidth));
    cos_rom(160) <= std_logic_vector(to_signed(-239,bitWidth));
    cos_rom(161) <= std_logic_vector(to_signed(-241,bitWidth));
    cos_rom(162) <= std_logic_vector(to_signed(-242,bitWidth));
    cos_rom(163) <= std_logic_vector(to_signed(-243,bitWidth));
    cos_rom(164) <= std_logic_vector(to_signed(-245,bitWidth));
    cos_rom(165) <= std_logic_vector(to_signed(-246,bitWidth));
    cos_rom(166) <= std_logic_vector(to_signed(-247,bitWidth));
    cos_rom(167) <= std_logic_vector(to_signed(-248,bitWidth));
    cos_rom(168) <= std_logic_vector(to_signed(-249,bitWidth));
    cos_rom(169) <= std_logic_vector(to_signed(-250,bitWidth));
    cos_rom(170) <= std_logic_vector(to_signed(-251,bitWidth));
    cos_rom(171) <= std_logic_vector(to_signed(-251,bitWidth));
    cos_rom(172) <= std_logic_vector(to_signed(-252,bitWidth));
    cos_rom(173) <= std_logic_vector(to_signed(-253,bitWidth));
    cos_rom(174) <= std_logic_vector(to_signed(-253,bitWidth));
    cos_rom(175) <= std_logic_vector(to_signed(-254,bitWidth));
    cos_rom(176) <= std_logic_vector(to_signed(-254,bitWidth));
    cos_rom(177) <= std_logic_vector(to_signed(-254,bitWidth));
    cos_rom(178) <= std_logic_vector(to_signed(-254,bitWidth));
    cos_rom(179) <= std_logic_vector(to_signed(-254,bitWidth));
    cos_rom(180) <= std_logic_vector(to_signed(-255,bitWidth));
    cos_rom(181) <= std_logic_vector(to_signed(-254,bitWidth));
    cos_rom(182) <= std_logic_vector(to_signed(-254,bitWidth));
    cos_rom(183) <= std_logic_vector(to_signed(-254,bitWidth));
    cos_rom(184) <= std_logic_vector(to_signed(-254,bitWidth));
    cos_rom(185) <= std_logic_vector(to_signed(-254,bitWidth));
    cos_rom(186) <= std_logic_vector(to_signed(-253,bitWidth));
    cos_rom(187) <= std_logic_vector(to_signed(-253,bitWidth));
    cos_rom(188) <= std_logic_vector(to_signed(-252,bitWidth));
    cos_rom(189) <= std_logic_vector(to_signed(-251,bitWidth));
    cos_rom(190) <= std_logic_vector(to_signed(-251,bitWidth));
    cos_rom(191) <= std_logic_vector(to_signed(-250,bitWidth));
    cos_rom(192) <= std_logic_vector(to_signed(-249,bitWidth));
    cos_rom(193) <= std_logic_vector(to_signed(-248,bitWidth));
    cos_rom(194) <= std_logic_vector(to_signed(-247,bitWidth));
    cos_rom(195) <= std_logic_vector(to_signed(-246,bitWidth));
    cos_rom(196) <= std_logic_vector(to_signed(-245,bitWidth));
    cos_rom(197) <= std_logic_vector(to_signed(-243,bitWidth));
    cos_rom(198) <= std_logic_vector(to_signed(-242,bitWidth));
    cos_rom(199) <= std_logic_vector(to_signed(-241,bitWidth));
    cos_rom(200) <= std_logic_vector(to_signed(-239,bitWidth));
    cos_rom(201) <= std_logic_vector(to_signed(-238,bitWidth));
    cos_rom(202) <= std_logic_vector(to_signed(-236,bitWidth));
    cos_rom(203) <= std_logic_vector(to_signed(-234,bitWidth));
    cos_rom(204) <= std_logic_vector(to_signed(-232,bitWidth));
    cos_rom(205) <= std_logic_vector(to_signed(-231,bitWidth));
    cos_rom(206) <= std_logic_vector(to_signed(-229,bitWidth));
    cos_rom(207) <= std_logic_vector(to_signed(-227,bitWidth));
    cos_rom(208) <= std_logic_vector(to_signed(-225,bitWidth));
    cos_rom(209) <= std_logic_vector(to_signed(-223,bitWidth));
    cos_rom(210) <= std_logic_vector(to_signed(-220,bitWidth));
    cos_rom(211) <= std_logic_vector(to_signed(-218,bitWidth));
    cos_rom(212) <= std_logic_vector(to_signed(-216,bitWidth));
    cos_rom(213) <= std_logic_vector(to_signed(-213,bitWidth));
    cos_rom(214) <= std_logic_vector(to_signed(-211,bitWidth));
    cos_rom(215) <= std_logic_vector(to_signed(-208,bitWidth));
    cos_rom(216) <= std_logic_vector(to_signed(-206,bitWidth));
    cos_rom(217) <= std_logic_vector(to_signed(-203,bitWidth));
    cos_rom(218) <= std_logic_vector(to_signed(-200,bitWidth));
    cos_rom(219) <= std_logic_vector(to_signed(-198,bitWidth));
    cos_rom(220) <= std_logic_vector(to_signed(-195,bitWidth));
    cos_rom(221) <= std_logic_vector(to_signed(-192,bitWidth));
    cos_rom(222) <= std_logic_vector(to_signed(-189,bitWidth));
    cos_rom(223) <= std_logic_vector(to_signed(-186,bitWidth));
    cos_rom(224) <= std_logic_vector(to_signed(-183,bitWidth));
    cos_rom(225) <= std_logic_vector(to_signed(-180,bitWidth));
    cos_rom(226) <= std_logic_vector(to_signed(-177,bitWidth));
    cos_rom(227) <= std_logic_vector(to_signed(-173,bitWidth));
    cos_rom(228) <= std_logic_vector(to_signed(-170,bitWidth));
    cos_rom(229) <= std_logic_vector(to_signed(-167,bitWidth));
    cos_rom(230) <= std_logic_vector(to_signed(-163,bitWidth));
    cos_rom(231) <= std_logic_vector(to_signed(-160,bitWidth));
    cos_rom(232) <= std_logic_vector(to_signed(-156,bitWidth));
    cos_rom(233) <= std_logic_vector(to_signed(-153,bitWidth));
    cos_rom(234) <= std_logic_vector(to_signed(-149,bitWidth));
    cos_rom(235) <= std_logic_vector(to_signed(-146,bitWidth));
    cos_rom(236) <= std_logic_vector(to_signed(-142,bitWidth));
    cos_rom(237) <= std_logic_vector(to_signed(-138,bitWidth));
    cos_rom(238) <= std_logic_vector(to_signed(-135,bitWidth));
    cos_rom(239) <= std_logic_vector(to_signed(-131,bitWidth));
    cos_rom(240) <= std_logic_vector(to_signed(-127,bitWidth));
    cos_rom(241) <= std_logic_vector(to_signed(-123,bitWidth));
    cos_rom(242) <= std_logic_vector(to_signed(-119,bitWidth));
    cos_rom(243) <= std_logic_vector(to_signed(-115,bitWidth));
    cos_rom(244) <= std_logic_vector(to_signed(-111,bitWidth));
    cos_rom(245) <= std_logic_vector(to_signed(-107,bitWidth));
    cos_rom(246) <= std_logic_vector(to_signed(-103,bitWidth));
    cos_rom(247) <= std_logic_vector(to_signed(-99,bitWidth));
    cos_rom(248) <= std_logic_vector(to_signed(-95,bitWidth));
    cos_rom(249) <= std_logic_vector(to_signed(-91,bitWidth));
    cos_rom(250) <= std_logic_vector(to_signed(-87,bitWidth));
    cos_rom(251) <= std_logic_vector(to_signed(-83,bitWidth));
    cos_rom(252) <= std_logic_vector(to_signed(-78,bitWidth));
    cos_rom(253) <= std_logic_vector(to_signed(-74,bitWidth));
    cos_rom(254) <= std_logic_vector(to_signed(-70,bitWidth));
    cos_rom(255) <= std_logic_vector(to_signed(-65,bitWidth));
    cos_rom(256) <= std_logic_vector(to_signed(-61,bitWidth));
    cos_rom(257) <= std_logic_vector(to_signed(-57,bitWidth));
    cos_rom(258) <= std_logic_vector(to_signed(-53,bitWidth));
    cos_rom(259) <= std_logic_vector(to_signed(-48,bitWidth));
    cos_rom(260) <= std_logic_vector(to_signed(-44,bitWidth));
    cos_rom(261) <= std_logic_vector(to_signed(-39,bitWidth));
    cos_rom(262) <= std_logic_vector(to_signed(-35,bitWidth));
    cos_rom(263) <= std_logic_vector(to_signed(-31,bitWidth));
    cos_rom(264) <= std_logic_vector(to_signed(-26,bitWidth));
    cos_rom(265) <= std_logic_vector(to_signed(-22,bitWidth));
    cos_rom(266) <= std_logic_vector(to_signed(-17,bitWidth));
    cos_rom(267) <= std_logic_vector(to_signed(-13,bitWidth));
    cos_rom(268) <= std_logic_vector(to_signed(-8,bitWidth));
    cos_rom(269) <= std_logic_vector(to_signed(-4,bitWidth));
    cos_rom(270) <= std_logic_vector(to_signed(0,bitWidth));
    cos_rom(271) <= std_logic_vector(to_signed(4,bitWidth));
    cos_rom(272) <= std_logic_vector(to_signed(8,bitWidth));
    cos_rom(273) <= std_logic_vector(to_signed(13,bitWidth));
    cos_rom(274) <= std_logic_vector(to_signed(17,bitWidth));
    cos_rom(275) <= std_logic_vector(to_signed(22,bitWidth));
    cos_rom(276) <= std_logic_vector(to_signed(26,bitWidth));
    cos_rom(277) <= std_logic_vector(to_signed(31,bitWidth));
    cos_rom(278) <= std_logic_vector(to_signed(35,bitWidth));
    cos_rom(279) <= std_logic_vector(to_signed(39,bitWidth));
    cos_rom(280) <= std_logic_vector(to_signed(44,bitWidth));
    cos_rom(281) <= std_logic_vector(to_signed(48,bitWidth));
    cos_rom(282) <= std_logic_vector(to_signed(53,bitWidth));
    cos_rom(283) <= std_logic_vector(to_signed(57,bitWidth));
    cos_rom(284) <= std_logic_vector(to_signed(61,bitWidth));
    cos_rom(285) <= std_logic_vector(to_signed(65,bitWidth));
    cos_rom(286) <= std_logic_vector(to_signed(70,bitWidth));
    cos_rom(287) <= std_logic_vector(to_signed(74,bitWidth));
    cos_rom(288) <= std_logic_vector(to_signed(78,bitWidth));
    cos_rom(289) <= std_logic_vector(to_signed(83,bitWidth));
    cos_rom(290) <= std_logic_vector(to_signed(87,bitWidth));
    cos_rom(291) <= std_logic_vector(to_signed(91,bitWidth));
    cos_rom(292) <= std_logic_vector(to_signed(95,bitWidth));
    cos_rom(293) <= std_logic_vector(to_signed(99,bitWidth));
    cos_rom(294) <= std_logic_vector(to_signed(103,bitWidth));
    cos_rom(295) <= std_logic_vector(to_signed(107,bitWidth));
    cos_rom(296) <= std_logic_vector(to_signed(111,bitWidth));
    cos_rom(297) <= std_logic_vector(to_signed(115,bitWidth));
    cos_rom(298) <= std_logic_vector(to_signed(119,bitWidth));
    cos_rom(299) <= std_logic_vector(to_signed(123,bitWidth));
    cos_rom(300) <= std_logic_vector(to_signed(127,bitWidth));
    cos_rom(301) <= std_logic_vector(to_signed(131,bitWidth));
    cos_rom(302) <= std_logic_vector(to_signed(135,bitWidth));
    cos_rom(303) <= std_logic_vector(to_signed(138,bitWidth));
    cos_rom(304) <= std_logic_vector(to_signed(142,bitWidth));
    cos_rom(305) <= std_logic_vector(to_signed(146,bitWidth));
    cos_rom(306) <= std_logic_vector(to_signed(149,bitWidth));
    cos_rom(307) <= std_logic_vector(to_signed(153,bitWidth));
    cos_rom(308) <= std_logic_vector(to_signed(156,bitWidth));
    cos_rom(309) <= std_logic_vector(to_signed(160,bitWidth));
    cos_rom(310) <= std_logic_vector(to_signed(163,bitWidth));
    cos_rom(311) <= std_logic_vector(to_signed(167,bitWidth));
    cos_rom(312) <= std_logic_vector(to_signed(170,bitWidth));
    cos_rom(313) <= std_logic_vector(to_signed(173,bitWidth));
    cos_rom(314) <= std_logic_vector(to_signed(177,bitWidth));
    cos_rom(315) <= std_logic_vector(to_signed(180,bitWidth));
    cos_rom(316) <= std_logic_vector(to_signed(183,bitWidth));
    cos_rom(317) <= std_logic_vector(to_signed(186,bitWidth));
    cos_rom(318) <= std_logic_vector(to_signed(189,bitWidth));
    cos_rom(319) <= std_logic_vector(to_signed(192,bitWidth));
    cos_rom(320) <= std_logic_vector(to_signed(195,bitWidth));
    cos_rom(321) <= std_logic_vector(to_signed(198,bitWidth));
    cos_rom(322) <= std_logic_vector(to_signed(200,bitWidth));
    cos_rom(323) <= std_logic_vector(to_signed(203,bitWidth));
    cos_rom(324) <= std_logic_vector(to_signed(206,bitWidth));
    cos_rom(325) <= std_logic_vector(to_signed(208,bitWidth));
    cos_rom(326) <= std_logic_vector(to_signed(211,bitWidth));
    cos_rom(327) <= std_logic_vector(to_signed(213,bitWidth));
    cos_rom(328) <= std_logic_vector(to_signed(216,bitWidth));
    cos_rom(329) <= std_logic_vector(to_signed(218,bitWidth));
    cos_rom(330) <= std_logic_vector(to_signed(220,bitWidth));
    cos_rom(331) <= std_logic_vector(to_signed(223,bitWidth));
    cos_rom(332) <= std_logic_vector(to_signed(225,bitWidth));
    cos_rom(333) <= std_logic_vector(to_signed(227,bitWidth));
    cos_rom(334) <= std_logic_vector(to_signed(229,bitWidth));
    cos_rom(335) <= std_logic_vector(to_signed(231,bitWidth));
    cos_rom(336) <= std_logic_vector(to_signed(232,bitWidth));
    cos_rom(337) <= std_logic_vector(to_signed(234,bitWidth));
    cos_rom(338) <= std_logic_vector(to_signed(236,bitWidth));
    cos_rom(339) <= std_logic_vector(to_signed(238,bitWidth));
    cos_rom(340) <= std_logic_vector(to_signed(239,bitWidth));
    cos_rom(341) <= std_logic_vector(to_signed(241,bitWidth));
    cos_rom(342) <= std_logic_vector(to_signed(242,bitWidth));
    cos_rom(343) <= std_logic_vector(to_signed(243,bitWidth));
    cos_rom(344) <= std_logic_vector(to_signed(245,bitWidth));
    cos_rom(345) <= std_logic_vector(to_signed(246,bitWidth));
    cos_rom(346) <= std_logic_vector(to_signed(247,bitWidth));
    cos_rom(347) <= std_logic_vector(to_signed(248,bitWidth));
    cos_rom(348) <= std_logic_vector(to_signed(249,bitWidth));
    cos_rom(349) <= std_logic_vector(to_signed(250,bitWidth));
    cos_rom(350) <= std_logic_vector(to_signed(251,bitWidth));
    cos_rom(351) <= std_logic_vector(to_signed(251,bitWidth));
    cos_rom(352) <= std_logic_vector(to_signed(252,bitWidth));
    cos_rom(353) <= std_logic_vector(to_signed(253,bitWidth));
    cos_rom(354) <= std_logic_vector(to_signed(253,bitWidth));
    cos_rom(355) <= std_logic_vector(to_signed(254,bitWidth));
    cos_rom(356) <= std_logic_vector(to_signed(254,bitWidth));
    cos_rom(357) <= std_logic_vector(to_signed(254,bitWidth));
    cos_rom(358) <= std_logic_vector(to_signed(254,bitWidth));
    cos_rom(359) <= std_logic_vector(to_signed(254,bitWidth));
    cos_rom(360) <= std_logic_vector(to_signed(255,bitWidth));
    report("trigo done");

end if;
end process;
end architecture;